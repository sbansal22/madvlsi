* SPICE3 file created from bias.ext - technology: sky130A


* Top level circuit bias

X0 a_600_1450# a_500_1420# a_n100_1450# a_n100_1450# sky130_fd_pr__nfet_01v8 ad=1.2e+13p pd=5.2e+07u as=4.2e+13p ps=1.82e+08u w=6e+06u l=500000u
X1 a_500_3170# a_500_3170# a_n100_1450# a_n100_1450# sky130_fd_pr__nfet_01v8 ad=6e+12p pd=2.6e+07u as=0p ps=0u w=6e+06u l=500000u
X2 a_600_4900# a_1100_4690# a_1100_4690# w_n140_4860# sky130_fd_pr__pfet_01v8 ad=1.2e+13p pd=5.2e+07u as=3e+12p ps=1.3e+07u w=6e+06u l=500000u
X3 w_n140_4860# w_n140_4860# w_n140_4860# w_n140_4860# sky130_fd_pr__pfet_01v8 ad=3.6e+13p pd=1.56e+08u as=0p ps=0u w=6e+06u l=500000u
X4 a_600_1450# a_500_1420# a_500_1420# a_n100_1450# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6e+12p ps=2.6e+07u w=6e+06u l=500000u
X5 w_n140_4860# a_140_6530# a_140_6530# w_n140_4860# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6e+12p ps=2.6e+07u w=6e+06u l=500000u
X6 a_400_3200# a_400_3200# a_600_4900# w_n140_4860# sky130_fd_pr__pfet_01v8 ad=6e+12p pd=2.6e+07u as=0p ps=0u w=6e+06u l=500000u
X7 a_400_3200# a_500_3170# a_n100_1450# a_n100_1450# sky130_fd_pr__nfet_01v8 ad=6e+12p pd=2.6e+07u as=0p ps=0u w=6e+06u l=500000u
X8 a_1100_4690# a_500_3170# a_n100_1450# a_n100_1450# sky130_fd_pr__nfet_01v8 ad=3e+12p pd=1.3e+07u as=0p ps=0u w=6e+06u l=500000u
X9 a_n100_1450# a_n100_1450# a_400_3200# a_n100_1450# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X10 a_n100_1450# a_n100_1450# a_n100_1450# a_n100_1450# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X11 a_800_6720# a_140_6530# w_n140_4860# w_n140_4860# sky130_fd_pr__pfet_01v8 ad=6e+12p pd=2.6e+07u as=0p ps=0u w=6e+06u l=500000u
X12 w_n140_4860# a_400_3200# a_600_4900# w_n140_4860# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X13 a_1100_4690# a_1100_4690# a_600_4900# w_n140_4860# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X14 a_n100_1450# a_500_3170# a_400_3200# a_n100_1450# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X15 w_n140_4860# w_n140_4860# w_n140_4860# w_n140_4860# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X16 w_n140_4860# a_140_6530# a_800_6720# w_n140_4860# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X17 a_140_6530# w_n140_4860# w_n140_4860# w_n140_4860# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X18 a_600_4900# a_400_3200# w_n140_4860# w_n140_4860# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X19 a_n100_1450# a_500_3170# a_500_3170# a_n100_1450# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X20 w_n140_4860# a_140_6530# a_500_1420# w_n140_4860# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3e+12p ps=1.3e+07u w=6e+06u l=500000u
X21 a_600_4900# a_400_3200# a_400_3200# w_n140_4860# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X22 a_n100_1450# a_n100_1450# a_n100_1450# a_n100_1450# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X23 a_400_3200# a_n100_1450# a_n100_1450# a_n100_1450# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X24 w_n140_4860# w_n140_4860# a_140_6530# w_n140_4860# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X25 a_600_1450# a_800_6720# a_800_6720# a_n100_1450# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3e+12p ps=1.3e+07u w=6e+06u l=500000u
X26 w_n140_4860# w_n140_4860# w_n140_4860# w_n140_4860# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X27 a_n100_1450# a_n100_1450# a_n100_1450# a_n100_1450# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X28 w_n140_4860# a_140_6530# a_500_3170# w_n140_4860# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6e+12p ps=2.6e+07u w=6e+06u l=500000u
X29 a_500_1420# a_500_1420# a_600_1450# a_n100_1450# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X30 a_500_1420# a_140_6530# w_n140_4860# w_n140_4860# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X31 a_n100_1450# a_n100_1450# a_n100_1450# a_n100_1450# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X32 a_140_6530# a_140_6530# w_n140_4860# w_n140_4860# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X33 a_n100_1450# a_500_1420# a_600_1450# a_n100_1450# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X34 a_500_3170# a_140_6530# w_n140_4860# w_n140_4860# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X35 a_800_6720# a_800_6720# a_600_1450# a_n100_1450# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X36 w_n140_4860# w_n140_4860# w_n140_4860# w_n140_4860# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X37 a_n100_1450# a_500_3170# a_1100_4690# a_n100_1450# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X38 a_n100_1450# a_n100_1450# a_n100_1450# a_n100_1450# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X39 a_n100_1450# a_n100_1450# a_n100_1450# a_n100_1450# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
.end

