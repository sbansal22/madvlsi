* SPICE3 file created from inverter-skinny.ext - technology: sky130A

.subckt inverter-skinny VP D VN CLK Dn
X0 Dn D VN VN sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X1 Dn D a_n340_1540# VP sky130_fd_pr__pfet_01v8 ad=9.025e+11p pd=5.7e+06u as=4.75e+11p ps=2.9e+06u w=950000u l=150000u
X2 Dn D a_n340_2000# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.75e+11p ps=2.9e+06u w=950000u l=150000u
.ends

