magic
tech sky130A
timestamp 1614289867
<< nmos >>
rect 25 1110 40 1205
rect 90 1110 105 1205
rect 155 1110 170 1205
rect 195 1110 210 1205
rect 25 785 40 880
rect 90 785 105 880
rect 155 785 170 880
rect 195 785 210 880
rect 25 520 40 620
rect 65 520 80 620
rect 130 520 145 620
rect 195 520 210 620
rect 25 170 40 270
rect 65 170 80 270
rect 130 170 145 270
rect 195 170 210 270
<< ndiff >>
rect -25 1190 25 1205
rect -25 1125 -10 1190
rect 10 1125 25 1190
rect -25 1110 25 1125
rect 40 1190 90 1205
rect 40 1125 55 1190
rect 75 1125 90 1190
rect 40 1110 90 1125
rect 105 1110 155 1205
rect 170 1110 195 1205
rect 210 1190 260 1205
rect 210 1125 225 1190
rect 245 1125 260 1190
rect 210 1110 260 1125
rect -25 865 25 880
rect -25 800 -10 865
rect 10 800 25 865
rect -25 785 25 800
rect 40 865 90 880
rect 40 800 55 865
rect 75 800 90 865
rect 40 785 90 800
rect 105 785 155 880
rect 170 785 195 880
rect 210 865 260 880
rect 210 800 225 865
rect 245 800 260 865
rect 210 785 260 800
rect -25 605 25 620
rect -25 535 -10 605
rect 10 535 25 605
rect -25 520 25 535
rect 40 520 65 620
rect 80 605 130 620
rect 80 535 95 605
rect 115 535 130 605
rect 80 520 130 535
rect 145 605 195 620
rect 145 535 160 605
rect 180 535 195 605
rect 145 520 195 535
rect 210 605 260 620
rect 210 535 225 605
rect 245 535 260 605
rect 210 520 260 535
rect -25 255 25 270
rect -25 185 -15 255
rect 10 185 25 255
rect -25 170 25 185
rect 40 170 65 270
rect 80 255 130 270
rect 80 185 95 255
rect 115 185 130 255
rect 80 170 130 185
rect 145 255 195 270
rect 145 185 160 255
rect 180 185 195 255
rect 145 170 195 185
rect 210 255 260 270
rect 210 185 225 255
rect 250 185 260 255
rect 210 170 260 185
<< ndiffc >>
rect -10 1125 10 1190
rect 55 1125 75 1190
rect 225 1125 245 1190
rect -10 800 10 865
rect 55 800 75 865
rect 225 800 245 865
rect -10 535 10 605
rect 95 535 115 605
rect 160 535 180 605
rect 225 535 245 605
rect -15 185 10 255
rect 95 185 115 255
rect 160 185 180 255
rect 225 185 250 255
<< psubdiff >>
rect -25 125 25 140
rect -25 55 -10 125
rect 10 55 25 125
rect -25 40 25 55
rect 210 125 260 140
rect 210 55 225 125
rect 245 55 260 125
rect 210 40 260 55
<< psubdiffcont >>
rect -10 55 10 125
rect 225 55 245 125
<< poly >>
rect 25 1205 40 1230
rect 90 1205 105 1230
rect 155 1205 170 1230
rect 195 1205 210 1230
rect 25 880 40 1110
rect 90 1055 105 1110
rect 155 1090 170 1110
rect 65 1045 105 1055
rect 65 1025 75 1045
rect 95 1025 105 1045
rect 65 1015 105 1025
rect 130 1075 170 1090
rect 65 980 105 990
rect 65 960 75 980
rect 95 960 105 980
rect 65 950 105 960
rect 90 880 105 950
rect 130 935 145 1075
rect 195 1050 210 1110
rect 170 1040 210 1050
rect 170 1020 180 1040
rect 200 1020 210 1040
rect 170 1010 210 1020
rect 130 920 170 935
rect 155 880 170 920
rect 195 925 250 935
rect 195 905 220 925
rect 240 905 250 925
rect 195 895 250 905
rect 195 880 210 895
rect 25 620 40 785
rect 90 775 105 785
rect 155 775 170 785
rect 65 760 105 775
rect 130 760 170 775
rect 65 620 80 760
rect 130 620 145 760
rect 195 620 210 785
rect 25 505 40 520
rect 0 490 40 505
rect 0 305 15 490
rect 65 465 80 520
rect 40 455 80 465
rect 40 435 50 455
rect 70 435 80 455
rect 40 425 80 435
rect 65 390 105 400
rect 65 370 75 390
rect 95 370 105 390
rect 65 360 105 370
rect 0 290 40 305
rect 25 270 40 290
rect 65 270 80 360
rect 130 270 145 520
rect 195 510 210 520
rect 170 495 210 510
rect 170 360 185 495
rect 210 460 250 470
rect 210 440 220 460
rect 240 440 250 460
rect 210 430 250 440
rect 170 350 210 360
rect 170 330 180 350
rect 200 330 210 350
rect 170 320 210 330
rect 235 295 250 430
rect 195 280 250 295
rect 195 270 210 280
rect 25 25 40 170
rect 65 155 80 170
rect 130 25 145 170
rect 195 155 210 170
rect 0 15 40 25
rect 0 -5 10 15
rect 30 -5 40 15
rect 0 -15 40 -5
rect 105 15 145 25
rect 105 -5 115 15
rect 135 -5 145 15
rect 105 -15 145 -5
<< polycont >>
rect 75 1025 95 1045
rect 75 960 95 980
rect 180 1020 200 1040
rect 220 905 240 925
rect 50 435 70 455
rect 75 370 95 390
rect 220 440 240 460
rect 180 330 200 350
rect 10 -5 30 15
rect 115 -5 135 15
<< locali >>
rect -25 1190 20 1200
rect -25 1125 -10 1190
rect 10 1125 20 1190
rect -25 1115 20 1125
rect 45 1190 85 1200
rect 45 1125 55 1190
rect 75 1125 85 1190
rect 45 1115 85 1125
rect 110 1115 150 1200
rect 215 1190 260 1200
rect 215 1125 225 1190
rect 245 1125 260 1190
rect 215 1115 260 1125
rect 65 1095 85 1115
rect 65 1075 145 1095
rect 65 1045 105 1055
rect 65 1035 75 1045
rect 25 1025 75 1035
rect 95 1025 105 1045
rect 25 1015 105 1025
rect 25 915 45 1015
rect 125 990 145 1075
rect 65 980 145 990
rect 65 960 75 980
rect 95 970 145 980
rect 170 1040 210 1050
rect 170 1020 180 1040
rect 200 1020 210 1040
rect 170 1010 210 1020
rect 95 960 105 970
rect 65 950 105 960
rect 25 895 65 915
rect 45 875 65 895
rect 170 875 190 1010
rect 230 935 250 1115
rect 210 925 250 935
rect 210 905 220 925
rect 240 905 250 925
rect 210 895 250 905
rect -25 865 20 875
rect -25 800 -10 865
rect 10 800 20 865
rect -25 790 20 800
rect 45 865 85 875
rect 45 800 55 865
rect 75 800 85 865
rect 45 790 85 800
rect 110 790 150 875
rect 170 865 260 875
rect 170 855 225 865
rect 215 800 225 855
rect 245 800 260 865
rect 65 615 85 790
rect 215 785 260 800
rect 215 780 235 785
rect 170 760 235 780
rect 170 615 190 760
rect -25 605 20 615
rect -25 535 -10 605
rect 10 535 20 605
rect 65 605 125 615
rect 65 590 95 605
rect -25 525 20 535
rect 85 535 95 590
rect 115 535 125 605
rect 85 525 125 535
rect 150 605 190 615
rect 150 535 160 605
rect 180 535 190 605
rect 150 525 190 535
rect 215 605 260 615
rect 215 535 225 605
rect 245 535 260 605
rect 215 525 260 535
rect 40 455 80 465
rect 40 445 50 455
rect 20 435 50 445
rect 70 435 80 455
rect 20 425 80 435
rect 20 335 40 425
rect 105 400 125 525
rect 170 470 190 525
rect 170 460 250 470
rect 170 450 220 460
rect 210 440 220 450
rect 240 440 250 460
rect 210 430 250 440
rect 65 390 125 400
rect 65 370 75 390
rect 95 380 125 390
rect 95 370 105 380
rect 65 360 105 370
rect 170 350 210 360
rect 20 315 105 335
rect 85 265 105 315
rect 170 330 180 350
rect 200 330 210 350
rect 170 320 210 330
rect 170 265 190 320
rect -25 255 20 265
rect -25 185 -15 255
rect 10 185 20 255
rect -25 175 20 185
rect 85 255 125 265
rect 85 185 95 255
rect 115 185 125 255
rect 85 175 125 185
rect 150 255 190 265
rect 150 185 160 255
rect 180 185 190 255
rect 150 175 190 185
rect 215 255 260 265
rect 215 185 225 255
rect 250 185 260 255
rect 215 175 260 185
rect -20 125 20 135
rect -20 55 -10 125
rect 10 55 20 125
rect -20 45 20 55
rect 215 125 255 135
rect 215 55 225 125
rect 245 55 255 125
rect 215 45 255 55
rect -25 15 260 25
rect -25 5 10 15
rect 0 -5 10 5
rect 30 5 115 15
rect 30 -5 40 5
rect 0 -15 40 -5
rect 105 -5 115 5
rect 135 5 260 15
rect 135 -5 145 5
rect 105 -15 145 -5
<< viali >>
rect -10 535 10 605
rect 225 535 245 605
rect -15 185 10 255
rect 225 185 250 255
rect -10 55 10 125
rect 225 55 245 125
<< metal1 >>
rect -25 605 20 620
rect -25 535 -10 605
rect 10 535 20 605
rect -25 255 20 535
rect -25 185 -15 255
rect 10 185 20 255
rect -25 140 20 185
rect 215 605 260 620
rect 215 535 225 605
rect 245 535 260 605
rect 215 255 260 535
rect 215 185 225 255
rect 250 185 260 255
rect 215 140 260 185
rect -25 125 260 140
rect -25 55 -10 125
rect 10 55 225 125
rect 245 55 260 125
rect -25 40 260 55
<< end >>
