magic
tech sky130A
timestamp 1613033220
<< nwell >>
rect -120 75 150 215
<< nmos >>
rect 0 -105 15 -5
rect 65 -105 80 -5
<< pmos >>
rect 0 95 15 195
rect 65 95 80 195
<< ndiff >>
rect -50 -20 0 -5
rect -50 -90 -35 -20
rect -15 -90 0 -20
rect -50 -105 0 -90
rect 15 -105 65 -5
rect 80 -20 130 -5
rect 80 -90 95 -20
rect 115 -90 130 -20
rect 80 -105 130 -90
<< pdiff >>
rect -50 180 0 195
rect -50 110 -35 180
rect -15 110 0 180
rect -50 95 0 110
rect 15 180 65 195
rect 15 110 30 180
rect 50 110 65 180
rect 15 95 65 110
rect 80 180 130 195
rect 80 110 95 180
rect 115 110 130 180
rect 80 95 130 110
<< ndiffc >>
rect -35 -90 -15 -20
rect 95 -90 115 -20
<< pdiffc >>
rect -35 110 -15 180
rect 30 110 50 180
rect 95 110 115 180
<< psubdiff >>
rect -100 -20 -50 -5
rect -100 -90 -85 -20
rect -65 -90 -50 -20
rect -100 -105 -50 -90
<< nsubdiff >>
rect -100 180 -50 195
rect -100 110 -85 180
rect -65 110 -50 180
rect -100 95 -50 110
<< psubdiffcont >>
rect -85 -90 -65 -20
<< nsubdiffcont >>
rect -85 110 -65 180
<< poly >>
rect 0 195 15 215
rect 65 195 80 215
rect 0 -5 15 95
rect 65 -5 80 95
rect 0 -120 15 -105
rect -25 -130 15 -120
rect -25 -150 -15 -130
rect 5 -150 15 -130
rect -25 -160 15 -150
rect 65 -185 80 -105
rect 40 -195 80 -185
rect 40 -215 50 -195
rect 70 -215 80 -195
rect 40 -225 80 -215
<< polycont >>
rect -15 -150 5 -130
rect 50 -215 70 -195
<< locali >>
rect -95 180 -5 190
rect -95 110 -85 180
rect -65 110 -35 180
rect -15 110 -5 180
rect -95 100 -5 110
rect 20 180 60 190
rect 20 110 30 180
rect 50 110 60 180
rect 20 100 60 110
rect 85 180 125 190
rect 85 110 95 180
rect 115 110 125 180
rect 85 100 125 110
rect -95 -20 -5 -10
rect -95 -90 -85 -20
rect -65 -90 -35 -20
rect -15 -90 -5 -20
rect -95 -100 -5 -90
rect 85 -20 125 -10
rect 85 -90 95 -20
rect 115 -90 125 -20
rect 85 -100 125 -90
rect 105 -120 125 -100
rect -120 -130 15 -120
rect -120 -140 -15 -130
rect -25 -150 -15 -140
rect 5 -150 15 -130
rect 105 -140 150 -120
rect -25 -160 15 -150
rect -120 -195 80 -185
rect -120 -205 50 -195
rect 40 -215 50 -205
rect 70 -215 80 -195
rect 40 -225 80 -215
<< viali >>
rect -85 110 -65 180
rect -35 110 -15 180
rect 95 110 115 180
rect -85 -90 -65 -20
rect -35 -90 -15 -20
<< metal1 >>
rect -120 180 150 190
rect -120 110 -85 180
rect -65 110 -35 180
rect -15 110 95 180
rect 115 110 150 180
rect -120 100 150 110
rect -120 -20 150 -10
rect -120 -90 -85 -20
rect -65 -90 -35 -20
rect -15 -90 150 -20
rect -120 -100 150 -90
<< labels >>
rlabel metal1 -120 -55 -120 -55 7 VN
port 5 w
rlabel metal1 -120 145 -120 145 7 VP
port 4 w
rlabel locali -120 -130 -120 -130 7 A
port 1 w
rlabel locali -120 -195 -120 -195 7 B
port 3 w
rlabel locali 150 -130 150 -130 3 Y
port 2 e
<< end >>
