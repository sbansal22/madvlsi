magic
tech sky130A
timestamp 1614683277
<< nwell >>
rect -45 855 280 1440
<< nmos >>
rect 25 620 40 820
rect 65 620 80 820
rect 130 620 145 720
rect 195 620 210 720
rect 25 170 40 370
rect 65 170 80 370
rect 130 270 145 370
rect 195 270 210 370
<< pmos >>
rect 25 1200 40 1295
rect 90 1200 105 1295
rect 155 1200 170 1295
rect 195 1200 210 1295
rect 25 875 40 970
rect 90 875 105 970
rect 155 875 170 970
rect 195 875 210 970
<< ndiff >>
rect -25 705 25 820
rect -25 635 -10 705
rect 10 635 25 705
rect -25 620 25 635
rect 40 620 65 820
rect 80 720 105 820
rect 80 705 130 720
rect 80 635 95 705
rect 115 635 130 705
rect 80 620 130 635
rect 145 705 195 720
rect 145 635 160 705
rect 180 635 195 705
rect 145 620 195 635
rect 210 705 260 720
rect 210 635 225 705
rect 245 635 260 705
rect 210 620 260 635
rect -25 355 25 370
rect -25 285 -15 355
rect 10 285 25 355
rect -25 170 25 285
rect 40 170 65 370
rect 80 355 130 370
rect 80 285 95 355
rect 115 285 130 355
rect 80 270 130 285
rect 145 355 195 370
rect 145 285 160 355
rect 180 285 195 355
rect 145 270 195 285
rect 210 355 260 370
rect 210 285 225 355
rect 250 285 260 355
rect 210 270 260 285
rect 80 170 105 270
<< pdiff >>
rect -25 1280 25 1295
rect -25 1215 -10 1280
rect 10 1215 25 1280
rect -25 1200 25 1215
rect 40 1280 90 1295
rect 40 1215 55 1280
rect 75 1215 90 1280
rect 40 1200 90 1215
rect 105 1280 155 1295
rect 105 1215 120 1280
rect 140 1215 155 1280
rect 105 1200 155 1215
rect 170 1200 195 1295
rect 210 1280 260 1295
rect 210 1215 225 1280
rect 245 1215 260 1280
rect 210 1200 260 1215
rect -25 955 25 970
rect -25 890 -10 955
rect 10 890 25 955
rect -25 875 25 890
rect 40 955 90 970
rect 40 890 55 955
rect 75 890 90 955
rect 40 875 90 890
rect 105 955 155 970
rect 105 890 120 955
rect 140 890 155 955
rect 105 875 155 890
rect 170 875 195 970
rect 210 955 260 970
rect 210 890 225 955
rect 245 890 260 955
rect 210 875 260 890
<< ndiffc >>
rect -10 635 10 705
rect 95 635 115 705
rect 160 635 180 705
rect 225 635 245 705
rect -15 285 10 355
rect 95 285 115 355
rect 160 285 180 355
rect 225 285 250 355
<< pdiffc >>
rect -10 1215 10 1280
rect 55 1215 75 1280
rect 120 1215 140 1280
rect 225 1215 245 1280
rect -10 890 10 955
rect 55 890 75 955
rect 120 890 140 955
rect 225 890 245 955
<< psubdiff >>
rect -25 125 25 140
rect -25 55 -10 125
rect 10 55 25 125
rect -25 40 25 55
rect 210 125 260 140
rect 210 55 225 125
rect 245 55 260 125
rect 210 40 260 55
<< nsubdiff >>
rect 105 1405 155 1420
rect 105 1340 120 1405
rect 140 1340 155 1405
rect 105 1325 155 1340
<< psubdiffcont >>
rect -10 55 10 125
rect 225 55 245 125
<< nsubdiffcont >>
rect 120 1340 140 1405
<< poly >>
rect 25 1295 40 1310
rect 90 1295 105 1310
rect 155 1295 170 1310
rect 195 1295 210 1310
rect 25 970 40 1200
rect 90 1145 105 1200
rect 155 1180 170 1200
rect 65 1135 105 1145
rect 65 1115 75 1135
rect 95 1115 105 1135
rect 65 1105 105 1115
rect 130 1165 170 1180
rect 65 1070 105 1080
rect 65 1050 75 1070
rect 95 1050 105 1070
rect 65 1040 105 1050
rect 90 970 105 1040
rect 130 1025 145 1165
rect 195 1140 210 1200
rect 170 1130 210 1140
rect 170 1110 180 1130
rect 200 1110 210 1130
rect 170 1100 210 1110
rect 130 1010 170 1025
rect 155 970 170 1010
rect 195 1015 250 1025
rect 195 995 220 1015
rect 240 995 250 1015
rect 195 985 250 995
rect 195 970 210 985
rect 25 820 40 875
rect 90 865 105 875
rect 155 865 170 875
rect 65 850 105 865
rect 130 850 170 865
rect 65 820 80 850
rect 130 720 145 850
rect 195 720 210 875
rect 25 605 40 620
rect 0 590 40 605
rect 0 405 15 590
rect 65 565 80 620
rect 40 555 80 565
rect 40 535 50 555
rect 70 535 80 555
rect 40 525 80 535
rect 65 490 105 500
rect 65 470 75 490
rect 95 470 105 490
rect 65 460 105 470
rect 0 390 40 405
rect 25 370 40 390
rect 65 370 80 460
rect 130 370 145 620
rect 195 610 210 620
rect 170 595 210 610
rect 170 460 185 595
rect 210 560 250 570
rect 210 540 220 560
rect 240 540 250 560
rect 210 530 250 540
rect 170 450 210 460
rect 170 430 180 450
rect 200 430 210 450
rect 170 420 210 430
rect 235 395 250 530
rect 195 380 250 395
rect 195 370 210 380
rect 25 25 40 170
rect 65 155 80 170
rect 130 25 145 270
rect 195 255 210 270
rect 0 15 40 25
rect 0 -5 10 15
rect 30 -5 40 15
rect 0 -15 40 -5
rect 105 15 145 25
rect 105 -5 115 15
rect 135 -5 145 15
rect 105 -15 145 -5
<< polycont >>
rect 75 1115 95 1135
rect 75 1050 95 1070
rect 180 1110 200 1130
rect 220 995 240 1015
rect 50 535 70 555
rect 75 470 95 490
rect 220 540 240 560
rect 180 430 200 450
rect 10 -5 30 15
rect 115 -5 135 15
<< locali >>
rect 110 1405 150 1415
rect 110 1340 120 1405
rect 140 1340 150 1405
rect 110 1330 150 1340
rect -25 1280 20 1290
rect -25 1260 -10 1280
rect -45 1240 -10 1260
rect -25 1215 -10 1240
rect 10 1215 20 1280
rect -25 1205 20 1215
rect 45 1280 85 1290
rect 45 1215 55 1280
rect 75 1215 85 1280
rect 45 1205 85 1215
rect 110 1280 150 1290
rect 110 1215 120 1280
rect 140 1215 150 1280
rect 110 1205 150 1215
rect 215 1280 260 1290
rect 215 1215 225 1280
rect 245 1260 260 1280
rect 245 1240 280 1260
rect 245 1215 260 1240
rect 215 1205 260 1215
rect 65 1185 85 1205
rect 65 1165 145 1185
rect 65 1135 105 1145
rect 65 1125 75 1135
rect 25 1115 75 1125
rect 95 1115 105 1135
rect 25 1105 105 1115
rect 25 1005 45 1105
rect 125 1080 145 1165
rect 65 1070 145 1080
rect 65 1050 75 1070
rect 95 1060 145 1070
rect 170 1130 210 1140
rect 170 1110 180 1130
rect 200 1110 210 1130
rect 170 1100 210 1110
rect 95 1050 105 1060
rect 65 1040 105 1050
rect 25 985 65 1005
rect 45 965 65 985
rect 170 965 190 1100
rect 230 1025 250 1205
rect 210 1015 250 1025
rect 210 995 220 1015
rect 240 995 250 1015
rect 210 985 250 995
rect -25 955 20 965
rect -25 935 -10 955
rect -45 915 -10 935
rect -25 890 -10 915
rect 10 890 20 955
rect -25 880 20 890
rect 45 955 85 965
rect 45 890 55 955
rect 75 890 85 955
rect 45 880 85 890
rect 110 955 150 965
rect 110 890 120 955
rect 140 890 150 955
rect 170 955 260 965
rect 170 945 225 955
rect 110 880 150 890
rect 215 890 225 945
rect 245 935 260 955
rect 245 915 280 935
rect 245 890 260 915
rect 65 715 85 880
rect 215 875 260 890
rect 215 870 235 875
rect 170 850 235 870
rect 170 715 190 850
rect -25 705 20 715
rect -25 635 -10 705
rect 10 635 20 705
rect 65 705 125 715
rect 65 690 95 705
rect -25 625 20 635
rect 85 635 95 690
rect 115 635 125 705
rect 85 625 125 635
rect 150 705 190 715
rect 150 635 160 705
rect 180 635 190 705
rect 150 625 190 635
rect 215 705 260 715
rect 215 635 225 705
rect 245 635 260 705
rect 215 625 260 635
rect 40 555 80 565
rect 40 545 50 555
rect 20 535 50 545
rect 70 535 80 555
rect 20 525 80 535
rect 20 435 40 525
rect 105 500 125 625
rect 170 570 190 625
rect 170 560 250 570
rect 170 550 220 560
rect 210 540 220 550
rect 240 540 250 560
rect 210 530 250 540
rect 65 490 125 500
rect 65 470 75 490
rect 95 480 125 490
rect 95 470 105 480
rect 65 460 105 470
rect 170 450 210 460
rect 20 415 105 435
rect 85 365 105 415
rect 170 430 180 450
rect 200 430 210 450
rect 170 420 210 430
rect 170 365 190 420
rect -25 355 20 365
rect -25 285 -15 355
rect 10 285 20 355
rect -25 275 20 285
rect 85 355 125 365
rect 85 285 95 355
rect 115 285 125 355
rect 85 275 125 285
rect 150 355 190 365
rect 150 285 160 355
rect 180 285 190 355
rect 150 275 190 285
rect 215 355 260 365
rect 215 285 225 355
rect 250 285 260 355
rect 215 275 260 285
rect -20 125 20 135
rect -20 55 -10 125
rect 10 55 20 125
rect -20 45 20 55
rect 215 125 255 135
rect 215 55 225 125
rect 245 55 255 125
rect 215 45 255 55
rect -45 15 280 25
rect -45 5 10 15
rect 0 -5 10 5
rect 30 5 115 15
rect 30 -5 40 5
rect 0 -15 40 -5
rect 105 -5 115 5
rect 135 5 280 15
rect 135 -5 145 5
rect 105 -15 145 -5
<< viali >>
rect 120 1340 140 1405
rect 120 1215 140 1280
rect 120 890 140 955
rect -10 635 10 705
rect 225 635 245 705
rect -15 285 10 355
rect 225 285 250 355
rect -10 55 10 125
rect 225 55 245 125
<< metal1 >>
rect -45 1405 280 1420
rect -45 1340 120 1405
rect 140 1340 280 1405
rect -45 1325 280 1340
rect 110 1280 150 1325
rect 110 1215 120 1280
rect 140 1215 150 1280
rect 110 955 150 1215
rect 110 890 120 955
rect 140 890 150 955
rect 110 880 150 890
rect -25 705 20 720
rect -25 635 -10 705
rect 10 635 20 705
rect -25 355 20 635
rect -25 285 -15 355
rect 10 285 20 355
rect -25 255 20 285
rect 215 705 260 720
rect 215 635 225 705
rect 245 635 260 705
rect 215 355 260 635
rect 215 285 225 355
rect 250 285 260 355
rect 215 255 260 285
rect -25 140 20 155
rect 215 140 260 155
rect -45 125 280 140
rect -45 55 -10 125
rect 10 55 225 125
rect 245 55 280 125
rect -45 40 280 55
<< labels >>
rlabel metal1 -45 90 -45 90 7 VN
port 4 w
rlabel locali -45 15 -45 15 7 CLK
port 5 w
rlabel locali 280 1250 280 1250 3 Qn
port 7 e
rlabel locali 280 925 280 925 3 Q
port 6 e
rlabel locali -45 925 -45 925 7 D
port 3 w
rlabel locali -45 1250 -45 1250 7 Dn
port 2 w
rlabel metal1 -45 1370 -45 1370 7 VP
port 1 w
<< end >>
