magic
tech sky130A
timestamp 1614290182
<< nmos >>
rect 25 1000 40 1095
rect 90 1000 105 1095
rect 155 1000 170 1095
rect 195 1000 210 1095
rect 25 675 40 770
rect 90 675 105 770
rect 155 675 170 770
rect 195 675 210 770
rect 25 520 40 620
rect 65 520 80 620
rect 130 520 145 620
rect 195 520 210 620
rect 25 170 40 270
rect 65 170 80 270
rect 130 170 145 270
rect 195 170 210 270
<< ndiff >>
rect -25 1080 25 1095
rect -25 1015 -10 1080
rect 10 1015 25 1080
rect -25 1000 25 1015
rect 40 1080 90 1095
rect 40 1015 55 1080
rect 75 1015 90 1080
rect 40 1000 90 1015
rect 105 1000 155 1095
rect 170 1000 195 1095
rect 210 1080 260 1095
rect 210 1015 225 1080
rect 245 1015 260 1080
rect 210 1000 260 1015
rect -25 755 25 770
rect -25 690 -10 755
rect 10 690 25 755
rect -25 675 25 690
rect 40 755 90 770
rect 40 690 55 755
rect 75 690 90 755
rect 40 675 90 690
rect 105 675 155 770
rect 170 675 195 770
rect 210 755 260 770
rect 210 690 225 755
rect 245 690 260 755
rect 210 675 260 690
rect -25 605 25 620
rect -25 535 -10 605
rect 10 535 25 605
rect -25 520 25 535
rect 40 520 65 620
rect 80 605 130 620
rect 80 535 95 605
rect 115 535 130 605
rect 80 520 130 535
rect 145 605 195 620
rect 145 535 160 605
rect 180 535 195 605
rect 145 520 195 535
rect 210 605 260 620
rect 210 535 225 605
rect 245 535 260 605
rect 210 520 260 535
rect -25 255 25 270
rect -25 185 -15 255
rect 10 185 25 255
rect -25 170 25 185
rect 40 170 65 270
rect 80 255 130 270
rect 80 185 95 255
rect 115 185 130 255
rect 80 170 130 185
rect 145 255 195 270
rect 145 185 160 255
rect 180 185 195 255
rect 145 170 195 185
rect 210 255 260 270
rect 210 185 225 255
rect 250 185 260 255
rect 210 170 260 185
<< ndiffc >>
rect -10 1015 10 1080
rect 55 1015 75 1080
rect 225 1015 245 1080
rect -10 690 10 755
rect 55 690 75 755
rect 225 690 245 755
rect -10 535 10 605
rect 95 535 115 605
rect 160 535 180 605
rect 225 535 245 605
rect -15 185 10 255
rect 95 185 115 255
rect 160 185 180 255
rect 225 185 250 255
<< psubdiff >>
rect -25 125 25 140
rect -25 55 -10 125
rect 10 55 25 125
rect -25 40 25 55
rect 210 125 260 140
rect 210 55 225 125
rect 245 55 260 125
rect 210 40 260 55
<< psubdiffcont >>
rect -10 55 10 125
rect 225 55 245 125
<< poly >>
rect 25 1095 40 1110
rect 90 1095 105 1110
rect 155 1095 170 1110
rect 195 1095 210 1110
rect 25 770 40 1000
rect 90 945 105 1000
rect 155 980 170 1000
rect 65 935 105 945
rect 65 915 75 935
rect 95 915 105 935
rect 65 905 105 915
rect 130 965 170 980
rect 65 870 105 880
rect 65 850 75 870
rect 95 850 105 870
rect 65 840 105 850
rect 90 770 105 840
rect 130 825 145 965
rect 195 940 210 1000
rect 170 930 210 940
rect 170 910 180 930
rect 200 910 210 930
rect 170 900 210 910
rect 130 810 170 825
rect 155 770 170 810
rect 195 815 250 825
rect 195 795 220 815
rect 240 795 250 815
rect 195 785 250 795
rect 195 770 210 785
rect 25 620 40 675
rect 90 665 105 675
rect 155 665 170 675
rect 65 650 105 665
rect 130 650 170 665
rect 65 620 80 650
rect 130 620 145 650
rect 195 620 210 675
rect 25 505 40 520
rect 0 490 40 505
rect 0 305 15 490
rect 65 465 80 520
rect 40 455 80 465
rect 40 435 50 455
rect 70 435 80 455
rect 40 425 80 435
rect 65 390 105 400
rect 65 370 75 390
rect 95 370 105 390
rect 65 360 105 370
rect 0 290 40 305
rect 25 270 40 290
rect 65 270 80 360
rect 130 270 145 520
rect 195 510 210 520
rect 170 495 210 510
rect 170 360 185 495
rect 210 460 250 470
rect 210 440 220 460
rect 240 440 250 460
rect 210 430 250 440
rect 170 350 210 360
rect 170 330 180 350
rect 200 330 210 350
rect 170 320 210 330
rect 235 295 250 430
rect 195 280 250 295
rect 195 270 210 280
rect 25 25 40 170
rect 65 155 80 170
rect 130 25 145 170
rect 195 155 210 170
rect 0 15 40 25
rect 0 -5 10 15
rect 30 -5 40 15
rect 0 -15 40 -5
rect 105 15 145 25
rect 105 -5 115 15
rect 135 -5 145 15
rect 105 -15 145 -5
<< polycont >>
rect 75 915 95 935
rect 75 850 95 870
rect 180 910 200 930
rect 220 795 240 815
rect 50 435 70 455
rect 75 370 95 390
rect 220 440 240 460
rect 180 330 200 350
rect 10 -5 30 15
rect 115 -5 135 15
<< locali >>
rect -25 1080 20 1090
rect -25 1015 -10 1080
rect 10 1015 20 1080
rect -25 1005 20 1015
rect 45 1080 85 1090
rect 45 1015 55 1080
rect 75 1015 85 1080
rect 45 1005 85 1015
rect 110 1005 150 1090
rect 215 1080 260 1090
rect 215 1015 225 1080
rect 245 1015 260 1080
rect 215 1005 260 1015
rect 65 985 85 1005
rect 65 965 145 985
rect 65 935 105 945
rect 65 925 75 935
rect 25 915 75 925
rect 95 915 105 935
rect 25 905 105 915
rect 25 805 45 905
rect 125 880 145 965
rect 65 870 145 880
rect 65 850 75 870
rect 95 860 145 870
rect 170 930 210 940
rect 170 910 180 930
rect 200 910 210 930
rect 170 900 210 910
rect 95 850 105 860
rect 65 840 105 850
rect 25 785 65 805
rect 45 765 65 785
rect 170 765 190 900
rect 230 825 250 1005
rect 210 815 250 825
rect 210 795 220 815
rect 240 795 250 815
rect 210 785 250 795
rect -25 755 20 765
rect -25 690 -10 755
rect 10 690 20 755
rect -25 680 20 690
rect 45 755 85 765
rect 45 690 55 755
rect 75 690 85 755
rect 45 680 85 690
rect 110 680 150 765
rect 170 755 260 765
rect 170 745 225 755
rect 215 690 225 745
rect 245 690 260 755
rect 65 615 85 680
rect 215 675 260 690
rect 215 670 235 675
rect 170 650 235 670
rect 170 615 190 650
rect -25 605 20 615
rect -25 535 -10 605
rect 10 535 20 605
rect 65 605 125 615
rect 65 590 95 605
rect -25 525 20 535
rect 85 535 95 590
rect 115 535 125 605
rect 85 525 125 535
rect 150 605 190 615
rect 150 535 160 605
rect 180 535 190 605
rect 150 525 190 535
rect 215 605 260 615
rect 215 535 225 605
rect 245 535 260 605
rect 215 525 260 535
rect 40 455 80 465
rect 40 445 50 455
rect 20 435 50 445
rect 70 435 80 455
rect 20 425 80 435
rect 20 335 40 425
rect 105 400 125 525
rect 170 470 190 525
rect 170 460 250 470
rect 170 450 220 460
rect 210 440 220 450
rect 240 440 250 460
rect 210 430 250 440
rect 65 390 125 400
rect 65 370 75 390
rect 95 380 125 390
rect 95 370 105 380
rect 65 360 105 370
rect 170 350 210 360
rect 20 315 105 335
rect 85 265 105 315
rect 170 330 180 350
rect 200 330 210 350
rect 170 320 210 330
rect 170 265 190 320
rect -25 255 20 265
rect -25 185 -15 255
rect 10 185 20 255
rect -25 175 20 185
rect 85 255 125 265
rect 85 185 95 255
rect 115 185 125 255
rect 85 175 125 185
rect 150 255 190 265
rect 150 185 160 255
rect 180 185 190 255
rect 150 175 190 185
rect 215 255 260 265
rect 215 185 225 255
rect 250 185 260 255
rect 215 175 260 185
rect -20 125 20 135
rect -20 55 -10 125
rect 10 55 20 125
rect -20 45 20 55
rect 215 125 255 135
rect 215 55 225 125
rect 245 55 255 125
rect 215 45 255 55
rect -25 15 260 25
rect -25 5 10 15
rect 0 -5 10 5
rect 30 5 115 15
rect 30 -5 40 5
rect 0 -15 40 -5
rect 105 -5 115 5
rect 135 5 260 15
rect 135 -5 145 5
rect 105 -15 145 -5
<< viali >>
rect -10 535 10 605
rect 225 535 245 605
rect -15 185 10 255
rect 225 185 250 255
rect -10 55 10 125
rect 225 55 245 125
<< metal1 >>
rect -25 1125 260 1220
rect 110 680 150 1125
rect -25 605 20 620
rect -25 535 -10 605
rect 10 535 20 605
rect -25 255 20 535
rect -25 185 -15 255
rect 10 185 20 255
rect -25 140 20 185
rect 215 605 260 620
rect 215 535 225 605
rect 245 535 260 605
rect 215 255 260 535
rect 215 185 225 255
rect 250 185 260 255
rect 215 140 260 185
rect -25 125 260 140
rect -25 55 -10 125
rect 10 55 225 125
rect 245 55 260 125
rect -25 40 260 55
<< end >>
