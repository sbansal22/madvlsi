magic
tech sky130A
timestamp 1615891844
<< nwell >>
rect -70 2430 1320 3980
<< nmos >>
rect 50 1600 100 2200
rect 150 1600 200 2200
rect 250 1600 300 2200
rect 350 1600 400 2200
rect 550 1600 600 2200
rect 650 1600 700 2200
rect 850 1600 900 2200
rect 950 1600 1000 2200
rect 1050 1600 1100 2200
rect 1150 1600 1200 2200
rect 50 725 100 1325
rect 150 725 200 1325
rect 250 725 300 1325
rect 350 725 400 1325
rect 550 725 600 1325
rect 650 725 700 1325
rect 850 725 900 1325
rect 950 725 1000 1325
rect 1050 725 1100 1325
rect 1150 725 1200 1325
<< pmos >>
rect 50 3360 100 3960
rect 150 3360 200 3960
rect 250 3360 300 3960
rect 450 3360 500 3960
rect 550 3360 600 3960
rect 650 3360 700 3960
rect 750 3360 800 3960
rect 950 3360 1000 3960
rect 1050 3360 1100 3960
rect 1150 3360 1200 3960
rect 50 2450 100 3050
rect 150 2450 200 3050
rect 250 2450 300 3050
rect 350 2450 400 3050
rect 550 2450 600 3050
rect 650 2450 700 3050
rect 850 2450 900 3050
rect 950 2450 1000 3050
rect 1050 2450 1100 3050
rect 1150 2450 1200 3050
<< ndiff >>
rect 0 2185 50 2200
rect 0 1615 15 2185
rect 35 1615 50 2185
rect 0 1600 50 1615
rect 100 2185 150 2200
rect 100 1615 115 2185
rect 135 1615 150 2185
rect 100 1600 150 1615
rect 200 2185 250 2200
rect 200 1615 215 2185
rect 235 1615 250 2185
rect 200 1600 250 1615
rect 300 2185 350 2200
rect 300 1615 315 2185
rect 335 1615 350 2185
rect 300 1600 350 1615
rect 400 2185 450 2200
rect 400 1615 415 2185
rect 435 1615 450 2185
rect 400 1600 450 1615
rect 500 2185 550 2200
rect 500 1615 515 2185
rect 535 1615 550 2185
rect 500 1600 550 1615
rect 600 2185 650 2200
rect 600 1615 615 2185
rect 635 1615 650 2185
rect 600 1600 650 1615
rect 700 2185 750 2200
rect 700 1615 715 2185
rect 735 1615 750 2185
rect 700 1600 750 1615
rect 800 2185 850 2200
rect 800 1615 815 2185
rect 835 1615 850 2185
rect 800 1600 850 1615
rect 900 2185 950 2200
rect 900 1615 915 2185
rect 935 1615 950 2185
rect 900 1600 950 1615
rect 1000 2185 1050 2200
rect 1000 1615 1015 2185
rect 1035 1615 1050 2185
rect 1000 1600 1050 1615
rect 1100 2185 1150 2200
rect 1100 1615 1115 2185
rect 1135 1615 1150 2185
rect 1100 1600 1150 1615
rect 1200 2185 1250 2200
rect 1200 1615 1215 2185
rect 1235 1615 1250 2185
rect 1200 1600 1250 1615
rect 0 1310 50 1325
rect 0 740 15 1310
rect 35 740 50 1310
rect 0 725 50 740
rect 100 1310 150 1325
rect 100 740 115 1310
rect 135 740 150 1310
rect 100 725 150 740
rect 200 1310 250 1325
rect 200 740 215 1310
rect 235 740 250 1310
rect 200 725 250 740
rect 300 1310 350 1325
rect 300 740 315 1310
rect 335 740 350 1310
rect 300 725 350 740
rect 400 1310 450 1325
rect 400 740 415 1310
rect 435 740 450 1310
rect 400 725 450 740
rect 500 1310 550 1325
rect 500 740 515 1310
rect 535 740 550 1310
rect 500 725 550 740
rect 600 1310 650 1325
rect 600 740 615 1310
rect 635 740 650 1310
rect 600 725 650 740
rect 700 1310 750 1325
rect 700 740 715 1310
rect 735 740 750 1310
rect 700 725 750 740
rect 800 1310 850 1325
rect 800 740 815 1310
rect 835 740 850 1310
rect 800 725 850 740
rect 900 1310 950 1325
rect 900 740 915 1310
rect 935 740 950 1310
rect 900 725 950 740
rect 1000 1310 1050 1325
rect 1000 740 1015 1310
rect 1035 740 1050 1310
rect 1000 725 1050 740
rect 1100 1310 1150 1325
rect 1100 740 1115 1310
rect 1135 740 1150 1310
rect 1100 725 1150 740
rect 1200 1310 1250 1325
rect 1200 740 1215 1310
rect 1235 740 1250 1310
rect 1200 725 1250 740
<< pdiff >>
rect 0 3945 50 3960
rect 0 3375 15 3945
rect 35 3375 50 3945
rect 0 3360 50 3375
rect 100 3945 150 3960
rect 100 3375 115 3945
rect 135 3375 150 3945
rect 100 3360 150 3375
rect 200 3945 250 3960
rect 200 3375 215 3945
rect 235 3375 250 3945
rect 200 3360 250 3375
rect 300 3945 350 3960
rect 300 3375 315 3945
rect 335 3375 350 3945
rect 300 3360 350 3375
rect 400 3945 450 3960
rect 400 3375 415 3945
rect 435 3375 450 3945
rect 400 3360 450 3375
rect 500 3945 550 3960
rect 500 3375 515 3945
rect 535 3375 550 3945
rect 500 3360 550 3375
rect 600 3945 650 3960
rect 600 3375 615 3945
rect 635 3375 650 3945
rect 600 3360 650 3375
rect 700 3945 750 3960
rect 700 3375 715 3945
rect 735 3375 750 3945
rect 700 3360 750 3375
rect 800 3945 850 3960
rect 800 3375 815 3945
rect 835 3375 850 3945
rect 800 3360 850 3375
rect 900 3945 950 3960
rect 900 3375 915 3945
rect 935 3375 950 3945
rect 900 3360 950 3375
rect 1000 3945 1050 3960
rect 1000 3375 1015 3945
rect 1035 3375 1050 3945
rect 1000 3360 1050 3375
rect 1100 3945 1150 3960
rect 1100 3375 1115 3945
rect 1135 3375 1150 3945
rect 1100 3360 1150 3375
rect 1200 3945 1250 3960
rect 1200 3375 1215 3945
rect 1235 3375 1250 3945
rect 1200 3360 1250 3375
rect 0 3035 50 3050
rect 0 2465 15 3035
rect 35 2465 50 3035
rect 0 2450 50 2465
rect 100 3035 150 3050
rect 100 2465 115 3035
rect 135 2465 150 3035
rect 100 2450 150 2465
rect 200 3035 250 3050
rect 200 2465 215 3035
rect 235 2465 250 3035
rect 200 2450 250 2465
rect 300 3035 350 3050
rect 300 2465 315 3035
rect 335 2465 350 3035
rect 300 2450 350 2465
rect 400 3035 450 3050
rect 400 2465 415 3035
rect 435 2465 450 3035
rect 400 2450 450 2465
rect 500 3035 550 3050
rect 500 2465 515 3035
rect 535 2465 550 3035
rect 500 2450 550 2465
rect 600 3035 650 3050
rect 600 2465 615 3035
rect 635 2465 650 3035
rect 600 2450 650 2465
rect 700 3035 750 3050
rect 700 2465 715 3035
rect 735 2465 750 3035
rect 700 2450 750 2465
rect 800 3035 850 3050
rect 800 2465 815 3035
rect 835 2465 850 3035
rect 800 2450 850 2465
rect 900 3035 950 3050
rect 900 2465 915 3035
rect 935 2465 950 3035
rect 900 2450 950 2465
rect 1000 3035 1050 3050
rect 1000 2465 1015 3035
rect 1035 2465 1050 3035
rect 1000 2450 1050 2465
rect 1100 3035 1150 3050
rect 1100 2465 1115 3035
rect 1135 2465 1150 3035
rect 1100 2450 1150 2465
rect 1200 3035 1250 3050
rect 1200 2465 1215 3035
rect 1235 2465 1250 3035
rect 1200 2450 1250 2465
<< ndiffc >>
rect 15 1615 35 2185
rect 115 1615 135 2185
rect 215 1615 235 2185
rect 315 1615 335 2185
rect 415 1615 435 2185
rect 515 1615 535 2185
rect 615 1615 635 2185
rect 715 1615 735 2185
rect 815 1615 835 2185
rect 915 1615 935 2185
rect 1015 1615 1035 2185
rect 1115 1615 1135 2185
rect 1215 1615 1235 2185
rect 15 740 35 1310
rect 115 740 135 1310
rect 215 740 235 1310
rect 315 740 335 1310
rect 415 740 435 1310
rect 515 740 535 1310
rect 615 740 635 1310
rect 715 740 735 1310
rect 815 740 835 1310
rect 915 740 935 1310
rect 1015 740 1035 1310
rect 1115 740 1135 1310
rect 1215 740 1235 1310
<< pdiffc >>
rect 15 3375 35 3945
rect 115 3375 135 3945
rect 215 3375 235 3945
rect 315 3375 335 3945
rect 415 3375 435 3945
rect 515 3375 535 3945
rect 615 3375 635 3945
rect 715 3375 735 3945
rect 815 3375 835 3945
rect 915 3375 935 3945
rect 1015 3375 1035 3945
rect 1115 3375 1135 3945
rect 1215 3375 1235 3945
rect 15 2465 35 3035
rect 115 2465 135 3035
rect 215 2465 235 3035
rect 315 2465 335 3035
rect 415 2465 435 3035
rect 515 2465 535 3035
rect 615 2465 635 3035
rect 715 2465 735 3035
rect 815 2465 835 3035
rect 915 2465 935 3035
rect 1015 2465 1035 3035
rect 1115 2465 1135 3035
rect 1215 2465 1235 3035
<< psubdiff >>
rect -50 2185 0 2200
rect -50 1615 -35 2185
rect -15 1615 0 2185
rect -50 1600 0 1615
rect 1250 2185 1300 2200
rect 1250 1615 1265 2185
rect 1285 1615 1300 2185
rect 1250 1600 1300 1615
rect -50 1310 0 1325
rect -50 740 -35 1310
rect -15 740 0 1310
rect -50 725 0 740
rect 1250 1310 1300 1325
rect 1250 740 1265 1310
rect 1285 740 1300 1310
rect 1250 725 1300 740
<< nsubdiff >>
rect -50 3945 0 3960
rect -50 3375 -35 3945
rect -15 3375 0 3945
rect -50 3360 0 3375
rect 1250 3945 1300 3960
rect 1250 3375 1265 3945
rect 1285 3375 1300 3945
rect 1250 3360 1300 3375
rect -50 3035 0 3050
rect -50 2465 -35 3035
rect -15 2465 0 3035
rect -50 2450 0 2465
rect 1250 3035 1300 3050
rect 1250 2465 1265 3035
rect 1285 2465 1300 3035
rect 1250 2450 1300 2465
<< psubdiffcont >>
rect -35 1615 -15 2185
rect 1265 1615 1285 2185
rect -35 740 -15 1310
rect 1265 740 1285 1310
<< nsubdiffcont >>
rect -35 3375 -15 3945
rect 1265 3375 1285 3945
rect -35 2465 -15 3035
rect 1265 2465 1285 3035
<< poly >>
rect 50 3960 100 3975
rect 150 3960 200 3975
rect 250 3960 300 3975
rect 450 3960 500 3975
rect 550 3960 600 3975
rect 650 3960 700 3975
rect 750 3960 800 3975
rect 950 3960 1000 3975
rect 1050 3960 1100 3975
rect 1150 3960 1200 3975
rect 50 3345 100 3360
rect 5 3335 100 3345
rect 5 3315 15 3335
rect 35 3330 100 3335
rect 150 3345 200 3360
rect 250 3345 300 3360
rect 450 3345 500 3360
rect 550 3345 600 3360
rect 650 3345 700 3360
rect 750 3345 800 3360
rect 950 3345 1000 3360
rect 1050 3345 1100 3360
rect 150 3330 1100 3345
rect 1150 3345 1200 3360
rect 1150 3335 1245 3345
rect 1150 3330 1215 3335
rect 35 3315 45 3330
rect 5 3305 45 3315
rect 150 3305 165 3330
rect 70 3295 165 3305
rect 70 3275 80 3295
rect 100 3290 165 3295
rect 1085 3305 1100 3330
rect 1205 3315 1215 3330
rect 1235 3315 1245 3335
rect 1205 3305 1245 3315
rect 1085 3295 1180 3305
rect 1085 3290 1150 3295
rect 100 3275 110 3290
rect 70 3265 110 3275
rect 1140 3275 1150 3290
rect 1170 3275 1180 3295
rect 1140 3265 1180 3275
rect 405 3135 845 3145
rect 405 3120 415 3135
rect 385 3115 415 3120
rect 435 3130 815 3135
rect 435 3115 445 3130
rect 385 3105 445 3115
rect 805 3115 815 3130
rect 835 3120 845 3135
rect 835 3115 865 3120
rect 805 3105 865 3115
rect 105 3095 145 3105
rect 105 3080 115 3095
rect 50 3075 115 3080
rect 135 3080 145 3095
rect 385 3080 400 3105
rect 605 3095 645 3105
rect 605 3080 615 3095
rect 135 3075 200 3080
rect 50 3065 200 3075
rect 50 3050 100 3065
rect 150 3050 200 3065
rect 250 3065 400 3080
rect 250 3050 300 3065
rect 350 3050 400 3065
rect 550 3075 615 3080
rect 635 3080 645 3095
rect 850 3080 865 3105
rect 1105 3095 1145 3105
rect 1105 3080 1115 3095
rect 635 3075 700 3080
rect 550 3065 700 3075
rect 550 3050 600 3065
rect 650 3050 700 3065
rect 850 3065 1000 3080
rect 850 3050 900 3065
rect 950 3050 1000 3065
rect 1050 3075 1115 3080
rect 1135 3080 1145 3095
rect 1135 3075 1200 3080
rect 1050 3065 1200 3075
rect 1050 3050 1100 3065
rect 1150 3050 1200 3065
rect 50 2435 100 2450
rect 150 2435 200 2450
rect 250 2335 300 2450
rect 350 2435 400 2450
rect 550 2375 600 2450
rect 650 2435 700 2450
rect 850 2435 900 2450
rect 950 2435 1000 2450
rect 1050 2435 1100 2450
rect 1150 2435 1200 2450
rect 550 2355 565 2375
rect 585 2355 600 2375
rect 550 2345 600 2355
rect 250 2315 265 2335
rect 285 2320 300 2335
rect 925 2335 965 2345
rect 925 2320 935 2335
rect 285 2315 935 2320
rect 955 2315 965 2335
rect 250 2305 965 2315
rect 985 2285 1210 2295
rect 985 2280 1180 2285
rect 405 2270 445 2280
rect 405 2255 415 2270
rect 105 2245 145 2255
rect 105 2230 115 2245
rect 50 2225 115 2230
rect 135 2230 145 2245
rect 385 2250 415 2255
rect 435 2255 445 2270
rect 805 2270 845 2280
rect 805 2255 815 2270
rect 435 2250 815 2255
rect 835 2255 845 2270
rect 835 2250 865 2255
rect 385 2240 865 2250
rect 385 2230 400 2240
rect 135 2225 200 2230
rect 50 2215 200 2225
rect 50 2200 100 2215
rect 150 2200 200 2215
rect 250 2215 400 2230
rect 250 2200 300 2215
rect 350 2200 400 2215
rect 550 2200 600 2240
rect 650 2200 700 2240
rect 850 2230 865 2240
rect 985 2230 1000 2280
rect 1170 2265 1180 2280
rect 1200 2265 1210 2285
rect 1170 2255 1210 2265
rect 1105 2245 1145 2255
rect 1105 2230 1115 2245
rect 850 2215 1000 2230
rect 850 2200 900 2215
rect 950 2200 1000 2215
rect 1050 2225 1115 2230
rect 1135 2230 1145 2245
rect 1135 2225 1200 2230
rect 1050 2215 1200 2225
rect 1050 2200 1100 2215
rect 1150 2200 1200 2215
rect 50 1585 100 1600
rect 150 1585 200 1600
rect 250 1585 300 1600
rect 350 1585 400 1600
rect 550 1585 600 1600
rect 650 1585 700 1600
rect 850 1585 900 1600
rect 950 1585 1000 1600
rect 1050 1585 1100 1600
rect 1150 1585 1200 1600
rect 550 1570 700 1585
rect 405 1395 445 1405
rect 405 1380 415 1395
rect 105 1370 145 1380
rect 105 1355 115 1370
rect 50 1350 115 1355
rect 135 1355 145 1370
rect 385 1375 415 1380
rect 435 1380 445 1395
rect 805 1395 845 1405
rect 805 1380 815 1395
rect 435 1375 815 1380
rect 835 1380 845 1395
rect 835 1375 865 1380
rect 385 1365 865 1375
rect 385 1355 400 1365
rect 135 1350 200 1355
rect 50 1340 200 1350
rect 50 1325 100 1340
rect 150 1325 200 1340
rect 250 1340 400 1355
rect 850 1355 865 1365
rect 1105 1370 1145 1380
rect 1105 1355 1115 1370
rect 850 1340 1000 1355
rect 250 1325 300 1340
rect 350 1325 400 1340
rect 550 1325 600 1340
rect 650 1325 700 1340
rect 850 1325 900 1340
rect 950 1325 1000 1340
rect 1050 1350 1115 1355
rect 1135 1355 1145 1370
rect 1135 1350 1200 1355
rect 1050 1340 1200 1350
rect 1050 1325 1100 1340
rect 1150 1325 1200 1340
rect 50 710 100 725
rect 150 710 200 725
rect 250 710 300 725
rect 350 710 400 725
rect 550 710 600 725
rect 650 710 700 725
rect 850 710 900 725
rect 950 710 1000 725
rect 1050 710 1100 725
rect 1150 710 1200 725
rect 550 700 700 710
rect 550 695 615 700
rect 605 680 615 695
rect 635 695 700 700
rect 635 680 645 695
rect 605 670 645 680
<< polycont >>
rect 15 3315 35 3335
rect 80 3275 100 3295
rect 1215 3315 1235 3335
rect 1150 3275 1170 3295
rect 415 3115 435 3135
rect 815 3115 835 3135
rect 115 3075 135 3095
rect 615 3075 635 3095
rect 1115 3075 1135 3095
rect 565 2355 585 2375
rect 265 2315 285 2335
rect 935 2315 955 2335
rect 115 2225 135 2245
rect 415 2250 435 2270
rect 815 2250 835 2270
rect 1180 2265 1200 2285
rect 1115 2225 1135 2245
rect 115 1350 135 1370
rect 415 1375 435 1395
rect 815 1375 835 1395
rect 1115 1350 1135 1370
rect 615 680 635 700
<< locali >>
rect 1105 3985 1300 4005
rect -45 3945 45 3955
rect -45 3375 -35 3945
rect -15 3375 15 3945
rect 35 3375 45 3945
rect -45 3365 45 3375
rect 5 3335 45 3365
rect 5 3315 15 3335
rect 35 3315 45 3335
rect 5 3305 45 3315
rect 105 3945 145 3955
rect 105 3375 115 3945
rect 135 3375 145 3945
rect 105 3305 145 3375
rect 205 3945 245 3955
rect 205 3375 215 3945
rect 235 3375 245 3945
rect 205 3360 245 3375
rect 305 3945 345 3955
rect 305 3375 315 3945
rect 335 3375 345 3945
rect 70 3295 145 3305
rect 70 3285 80 3295
rect -50 3275 80 3285
rect 100 3275 145 3295
rect -50 3265 145 3275
rect 305 3205 345 3375
rect 405 3945 445 3955
rect 405 3375 415 3945
rect 435 3375 445 3945
rect 405 3240 445 3375
rect 505 3945 545 3955
rect 505 3375 515 3945
rect 535 3375 545 3945
rect 505 3365 545 3375
rect 605 3945 645 3955
rect 605 3375 615 3945
rect 635 3375 645 3945
rect 605 3295 645 3375
rect 705 3945 745 3955
rect 705 3375 715 3945
rect 735 3375 745 3945
rect 705 3365 745 3375
rect 805 3945 845 3955
rect 805 3375 815 3945
rect 835 3375 845 3945
rect 605 3275 615 3295
rect 635 3275 645 3295
rect 605 3265 645 3275
rect 805 3250 845 3375
rect 805 3240 815 3250
rect 405 3230 815 3240
rect 835 3230 845 3250
rect 405 3220 845 3230
rect 905 3945 945 3955
rect 905 3375 915 3945
rect 935 3375 945 3945
rect 305 3185 315 3205
rect 335 3195 345 3205
rect 905 3195 945 3375
rect 1005 3945 1045 3955
rect 1005 3375 1015 3945
rect 1035 3375 1045 3945
rect 1005 3365 1045 3375
rect 1105 3945 1145 3985
rect 1105 3375 1115 3945
rect 1135 3375 1145 3945
rect 1105 3305 1145 3375
rect 1205 3945 1295 3955
rect 1205 3375 1215 3945
rect 1235 3375 1265 3945
rect 1285 3375 1295 3945
rect 1205 3365 1295 3375
rect 1205 3335 1245 3365
rect 1205 3315 1215 3335
rect 1235 3315 1245 3335
rect 1205 3305 1245 3315
rect 1105 3295 1180 3305
rect 1105 3275 1150 3295
rect 1170 3275 1180 3295
rect 1105 3265 1180 3275
rect 335 3185 945 3195
rect 305 3175 945 3185
rect 405 3135 445 3145
rect 405 3115 415 3135
rect 435 3115 445 3135
rect 105 3095 145 3105
rect 105 3085 115 3095
rect 5 3075 115 3085
rect 135 3075 145 3095
rect 5 3065 145 3075
rect 5 3045 45 3065
rect -45 3035 45 3045
rect -45 2465 -35 3035
rect -15 2465 15 3035
rect 35 2465 45 3035
rect -45 2455 45 2465
rect 105 3035 145 3065
rect 105 2465 115 3035
rect 135 2465 145 3035
rect 105 2455 145 2465
rect 205 3035 245 3045
rect 205 2465 215 3035
rect 235 2465 245 3035
rect 205 2455 245 2465
rect 305 3035 345 3045
rect 305 2465 315 3035
rect 335 2465 345 3035
rect 305 2430 345 2465
rect 405 3035 445 3115
rect 805 3135 845 3145
rect 805 3115 815 3135
rect 835 3115 845 3135
rect 605 3095 645 3105
rect 605 3075 615 3095
rect 635 3075 645 3095
rect 405 2465 415 3035
rect 435 2465 445 3035
rect 405 2455 445 2465
rect 505 3035 545 3045
rect 505 2465 515 3035
rect 535 2465 545 3035
rect 505 2430 545 2465
rect 605 3035 645 3075
rect 605 2465 615 3035
rect 635 2465 645 3035
rect 605 2455 645 2465
rect 705 3035 745 3045
rect 705 2465 715 3035
rect 735 2465 745 3035
rect 705 2430 745 2465
rect 805 3035 845 3115
rect 1105 3095 1145 3105
rect 1105 3075 1115 3095
rect 1135 3085 1145 3095
rect 1135 3075 1245 3085
rect 1105 3065 1245 3075
rect 805 2465 815 3035
rect 835 2465 845 3035
rect 805 2455 845 2465
rect 905 3035 945 3045
rect 905 2465 915 3035
rect 935 2465 945 3035
rect 905 2430 945 2465
rect 1005 3035 1045 3045
rect 1005 2465 1015 3035
rect 1035 2465 1045 3035
rect 1005 2455 1045 2465
rect 1105 3035 1145 3065
rect 1105 2465 1115 3035
rect 1135 2465 1145 3035
rect 1105 2455 1145 2465
rect 1205 3045 1245 3065
rect 1205 3035 1295 3045
rect 1205 2465 1215 3035
rect 1235 2465 1265 3035
rect 1285 2465 1295 3035
rect 1205 2455 1295 2465
rect 305 2410 945 2430
rect 405 2375 445 2385
rect 405 2355 415 2375
rect 435 2355 445 2375
rect 250 2335 300 2345
rect 250 2325 265 2335
rect 205 2315 265 2325
rect 285 2315 300 2335
rect 205 2305 300 2315
rect 105 2245 145 2255
rect 105 2235 115 2245
rect 5 2225 115 2235
rect 135 2225 145 2245
rect 5 2215 145 2225
rect 5 2195 45 2215
rect -45 2185 45 2195
rect -45 1615 -35 2185
rect -15 1615 15 2185
rect 35 1615 45 2185
rect -45 1605 45 1615
rect 105 2185 145 2215
rect 105 1615 115 2185
rect 135 1615 145 2185
rect 105 1605 145 1615
rect 205 2185 245 2305
rect 405 2270 445 2355
rect 550 2375 1300 2385
rect 550 2355 565 2375
rect 585 2365 1300 2375
rect 585 2355 645 2365
rect 550 2345 645 2355
rect 405 2250 415 2270
rect 435 2250 445 2270
rect 205 1615 215 2185
rect 235 1615 245 2185
rect 205 1605 245 1615
rect 305 2185 345 2195
rect 305 1615 315 2185
rect 335 1615 345 2185
rect 305 1605 345 1615
rect 405 2185 445 2250
rect 405 1615 415 2185
rect 435 1615 445 2185
rect 405 1605 445 1615
rect 505 2185 545 2195
rect 505 1615 515 2185
rect 535 1615 545 2185
rect 505 1575 545 1615
rect 605 2185 645 2345
rect 925 2335 965 2345
rect 925 2315 935 2335
rect 955 2325 965 2335
rect 955 2315 1045 2325
rect 925 2305 1045 2315
rect 805 2270 845 2280
rect 805 2250 815 2270
rect 835 2250 845 2270
rect 605 1615 615 2185
rect 635 1615 645 2185
rect 605 1605 645 1615
rect 705 2185 745 2195
rect 705 1615 715 2185
rect 735 1615 745 2185
rect 705 1575 745 1615
rect 805 2185 845 2250
rect 805 1615 815 2185
rect 835 1615 845 2185
rect 805 1605 845 1615
rect 905 2185 945 2195
rect 905 1615 915 2185
rect 935 1615 945 2185
rect 905 1605 945 1615
rect 1005 2185 1045 2305
rect 1170 2285 1300 2295
rect 1170 2265 1180 2285
rect 1200 2275 1300 2285
rect 1200 2265 1210 2275
rect 1170 2255 1210 2265
rect 1005 1615 1015 2185
rect 1035 1615 1045 2185
rect 1005 1605 1045 1615
rect 1105 2245 1145 2255
rect 1105 2225 1115 2245
rect 1135 2235 1145 2245
rect 1135 2225 1245 2235
rect 1105 2215 1245 2225
rect 1105 2185 1145 2215
rect 1105 1615 1115 2185
rect 1135 1615 1145 2185
rect 1105 1605 1145 1615
rect 1205 2195 1245 2215
rect 1205 2185 1295 2195
rect 1205 1615 1215 2185
rect 1235 1615 1265 2185
rect 1285 1615 1295 2185
rect 1205 1605 1295 1615
rect 505 1555 745 1575
rect 305 1485 945 1505
rect 105 1370 145 1380
rect 105 1360 115 1370
rect 5 1350 115 1360
rect 135 1350 145 1370
rect 5 1340 145 1350
rect 5 1320 45 1340
rect -45 1310 45 1320
rect -45 740 -35 1310
rect -15 740 15 1310
rect 35 740 45 1310
rect -45 730 45 740
rect 105 1310 145 1340
rect 105 740 115 1310
rect 135 740 145 1310
rect 105 730 145 740
rect 205 1310 245 1320
rect 205 740 215 1310
rect 235 740 245 1310
rect 205 730 245 740
rect 305 1310 345 1485
rect 305 740 315 1310
rect 335 740 345 1310
rect 305 730 345 740
rect 405 1455 445 1465
rect 405 1435 415 1455
rect 435 1435 445 1455
rect 405 1395 445 1435
rect 405 1375 415 1395
rect 435 1375 445 1395
rect 405 1310 445 1375
rect 405 740 415 1310
rect 435 740 445 1310
rect 405 730 445 740
rect 505 1310 545 1485
rect 505 740 515 1310
rect 535 740 545 1310
rect 505 730 545 740
rect 605 1455 645 1465
rect 605 1435 615 1455
rect 635 1435 645 1455
rect 605 1310 645 1435
rect 605 740 615 1310
rect 635 740 645 1310
rect 605 700 645 740
rect 705 1310 745 1485
rect 705 740 715 1310
rect 735 740 745 1310
rect 705 730 745 740
rect 805 1395 845 1405
rect 805 1375 815 1395
rect 835 1375 845 1395
rect 805 1310 845 1375
rect 805 740 815 1310
rect 835 740 845 1310
rect 805 730 845 740
rect 905 1310 945 1485
rect 1105 1370 1145 1380
rect 1105 1350 1115 1370
rect 1135 1360 1145 1370
rect 1135 1350 1245 1360
rect 1105 1340 1245 1350
rect 905 740 915 1310
rect 935 740 945 1310
rect 905 730 945 740
rect 1005 1310 1045 1320
rect 1005 740 1015 1310
rect 1035 740 1045 1310
rect 1005 730 1045 740
rect 1105 1310 1145 1340
rect 1105 740 1115 1310
rect 1135 740 1145 1310
rect 1105 730 1145 740
rect 1205 1320 1245 1340
rect 1205 1310 1295 1320
rect 1205 740 1215 1310
rect 1235 740 1265 1310
rect 1285 740 1295 1310
rect 1205 730 1295 740
rect 605 680 615 700
rect 635 680 1300 700
rect 605 670 645 680
<< viali >>
rect -35 3375 -15 3945
rect 15 3375 35 3945
rect 215 3375 235 3945
rect 515 3375 535 3945
rect 715 3375 735 3945
rect 615 3275 635 3295
rect 815 3230 835 3250
rect 315 3185 335 3205
rect 1015 3375 1035 3945
rect 1215 3375 1235 3945
rect 1265 3375 1285 3945
rect -35 2465 -15 3030
rect 15 2465 35 3030
rect 115 2465 135 3035
rect 215 2465 235 3035
rect 1015 2465 1035 3035
rect 1115 2465 1135 3035
rect 1215 2465 1235 3035
rect 1265 2465 1285 3035
rect 415 2355 435 2375
rect -35 1615 -15 2185
rect 15 1615 35 2185
rect 115 1615 135 2185
rect 315 1615 335 2185
rect 515 1615 535 2185
rect 915 1615 935 2185
rect 1115 1615 1135 2185
rect 1215 1615 1235 2185
rect 1265 1615 1285 2185
rect -35 740 -15 1310
rect 15 740 35 1310
rect 115 740 135 1310
rect 215 740 235 1310
rect 415 1435 435 1455
rect 615 1435 635 1455
rect 1015 740 1035 1310
rect 1115 740 1135 1310
rect 1215 740 1235 1310
rect 1265 740 1285 1310
<< metal1 >>
rect -50 3945 1300 3955
rect -50 3375 -35 3945
rect -15 3375 15 3945
rect 35 3375 215 3945
rect 235 3375 515 3945
rect 535 3375 715 3945
rect 735 3375 1015 3945
rect 1035 3375 1215 3945
rect 1235 3375 1265 3945
rect 1285 3375 1300 3945
rect -50 3360 1300 3375
rect -50 3035 250 3360
rect 605 3295 645 3305
rect 605 3275 615 3295
rect 635 3275 645 3295
rect -50 3030 115 3035
rect -50 2465 -35 3030
rect -15 2465 15 3030
rect 35 2465 115 3030
rect 135 2465 215 3035
rect 235 2465 250 3035
rect -50 2455 250 2465
rect 305 3205 345 3215
rect 305 3185 315 3205
rect 335 3185 345 3205
rect 305 2385 345 3185
rect 305 2375 445 2385
rect 305 2355 415 2375
rect 435 2355 445 2375
rect 305 2345 445 2355
rect -50 2185 550 2195
rect -50 1615 -35 2185
rect -15 1615 15 2185
rect 35 1615 115 2185
rect 135 1615 315 2185
rect 335 1615 515 2185
rect 535 1615 550 2185
rect -50 1600 550 1615
rect -50 1320 350 1600
rect 605 1530 645 3275
rect 405 1490 645 1530
rect 805 3250 845 3260
rect 805 3230 815 3250
rect 835 3230 845 3250
rect 405 1455 445 1490
rect 805 1465 845 3230
rect 1000 3035 1300 3360
rect 1000 2465 1015 3035
rect 1035 2465 1115 3035
rect 1135 2465 1215 3035
rect 1235 2465 1265 3035
rect 1285 2465 1300 3035
rect 1000 2455 1300 2465
rect 405 1435 415 1455
rect 435 1435 445 1455
rect 405 1425 445 1435
rect 605 1455 845 1465
rect 605 1435 615 1455
rect 635 1435 845 1455
rect 605 1425 845 1435
rect 900 2185 1300 2195
rect 900 1615 915 2185
rect 935 1615 1115 2185
rect 1135 1615 1215 2185
rect 1235 1615 1265 2185
rect 1285 1615 1300 2185
rect 900 1320 1300 1615
rect -50 1310 1300 1320
rect -50 740 -35 1310
rect -15 740 15 1310
rect 35 740 115 1310
rect 135 740 215 1310
rect 235 740 1015 1310
rect 1035 740 1115 1310
rect 1135 740 1215 1310
rect 1235 740 1265 1310
rect 1285 740 1300 1310
rect -50 730 1300 740
<< labels >>
rlabel metal1 -50 3660 -50 3660 7 VP
port 1 w
rlabel metal1 -50 3275 -50 3275 7 Vbp
port 2 w
rlabel metal1 -50 1900 -50 1900 7 VN
port 3 w
rlabel locali 1300 690 1300 690 3 Vcn
port 4 e
rlabel locali 1300 2285 1300 2285 3 Vbn
port 5 e
rlabel locali 1300 2375 1300 2375 3 Vcp
port 6 e
rlabel locali 1300 3995 1300 3995 3 Vbp
port 7 e
<< end >>
