magic
tech sky130A
timestamp 1615890655
<< nwell >>
rect -750 1245 440 2795
<< nmos >>
rect -630 -460 -580 140
rect -530 -460 -480 140
rect -430 -460 -380 140
rect -330 -460 -280 140
rect -230 -460 -180 140
rect -130 -460 -80 140
rect -30 -460 20 140
rect 70 -460 120 140
rect 170 -460 220 140
rect 270 -460 320 140
<< pmos >>
rect -630 2640 -580 2775
rect -530 2640 -480 2775
rect -430 2640 -380 2775
rect -330 2640 -280 2775
rect -230 2640 -180 2775
rect -130 2640 -80 2775
rect -30 2640 20 2775
rect 70 2640 120 2775
rect 170 2640 220 2775
rect 270 2640 320 2775
rect -630 2140 -580 2440
rect -530 2140 -480 2440
rect -430 2140 -380 2440
rect -330 2140 -280 2440
rect -230 2140 -180 2440
rect -130 2140 -80 2440
rect -30 2140 20 2440
rect 70 2140 120 2440
rect 170 2140 220 2440
rect 270 2140 320 2440
rect -630 1265 -580 1865
rect -530 1265 -480 1865
rect -430 1265 -380 1865
rect -330 1265 -280 1865
rect -230 1265 -180 1865
rect -130 1265 -80 1865
rect -30 1265 20 1865
rect 70 1265 120 1865
rect 170 1265 220 1865
rect 270 1265 320 1865
<< ndiff >>
rect -680 125 -630 140
rect -680 -445 -665 125
rect -645 -445 -630 125
rect -680 -460 -630 -445
rect -580 125 -530 140
rect -580 -445 -565 125
rect -545 -445 -530 125
rect -580 -460 -530 -445
rect -480 125 -430 140
rect -480 -445 -465 125
rect -445 -445 -430 125
rect -480 -460 -430 -445
rect -380 125 -330 140
rect -380 -445 -365 125
rect -345 -445 -330 125
rect -380 -460 -330 -445
rect -280 125 -230 140
rect -280 -445 -265 125
rect -245 -445 -230 125
rect -280 -460 -230 -445
rect -180 125 -130 140
rect -180 -445 -165 125
rect -145 -445 -130 125
rect -180 -460 -130 -445
rect -80 125 -30 140
rect -80 -445 -65 125
rect -45 -445 -30 125
rect -80 -460 -30 -445
rect 20 125 70 140
rect 20 -445 35 125
rect 55 -445 70 125
rect 20 -460 70 -445
rect 120 125 170 140
rect 120 -445 135 125
rect 155 -445 170 125
rect 120 -460 170 -445
rect 220 125 270 140
rect 220 -445 235 125
rect 255 -445 270 125
rect 220 -460 270 -445
rect 320 125 370 140
rect 320 -445 335 125
rect 355 -445 370 125
rect 320 -460 370 -445
<< pdiff >>
rect -680 2760 -630 2775
rect -680 2655 -665 2760
rect -645 2655 -630 2760
rect -680 2640 -630 2655
rect -580 2760 -530 2775
rect -580 2655 -565 2760
rect -545 2655 -530 2760
rect -580 2640 -530 2655
rect -480 2760 -430 2775
rect -480 2655 -465 2760
rect -445 2655 -430 2760
rect -480 2640 -430 2655
rect -380 2760 -330 2775
rect -380 2655 -365 2760
rect -345 2655 -330 2760
rect -380 2640 -330 2655
rect -280 2760 -230 2775
rect -280 2655 -265 2760
rect -245 2655 -230 2760
rect -280 2640 -230 2655
rect -180 2760 -130 2775
rect -180 2655 -165 2760
rect -145 2655 -130 2760
rect -180 2640 -130 2655
rect -80 2760 -30 2775
rect -80 2655 -65 2760
rect -45 2655 -30 2760
rect -80 2640 -30 2655
rect 20 2760 70 2775
rect 20 2655 35 2760
rect 55 2655 70 2760
rect 20 2640 70 2655
rect 120 2760 170 2775
rect 120 2655 135 2760
rect 155 2655 170 2760
rect 120 2640 170 2655
rect 220 2760 270 2775
rect 220 2655 235 2760
rect 255 2655 270 2760
rect 220 2640 270 2655
rect 320 2760 370 2775
rect 320 2655 335 2760
rect 355 2655 370 2760
rect 320 2640 370 2655
rect -680 2425 -630 2440
rect -680 2155 -665 2425
rect -645 2155 -630 2425
rect -680 2140 -630 2155
rect -580 2425 -530 2440
rect -580 2155 -565 2425
rect -545 2155 -530 2425
rect -580 2140 -530 2155
rect -480 2425 -430 2440
rect -480 2155 -465 2425
rect -445 2155 -430 2425
rect -480 2140 -430 2155
rect -380 2425 -330 2440
rect -380 2155 -365 2425
rect -345 2155 -330 2425
rect -380 2140 -330 2155
rect -280 2425 -230 2440
rect -280 2155 -265 2425
rect -245 2155 -230 2425
rect -280 2140 -230 2155
rect -180 2425 -130 2440
rect -180 2155 -165 2425
rect -145 2155 -130 2425
rect -180 2140 -130 2155
rect -80 2425 -30 2440
rect -80 2155 -65 2425
rect -45 2155 -30 2425
rect -80 2140 -30 2155
rect 20 2425 70 2440
rect 20 2155 35 2425
rect 55 2155 70 2425
rect 20 2140 70 2155
rect 120 2425 170 2440
rect 120 2155 135 2425
rect 155 2155 170 2425
rect 120 2140 170 2155
rect 220 2425 270 2440
rect 220 2155 235 2425
rect 255 2155 270 2425
rect 220 2140 270 2155
rect 320 2425 370 2440
rect 320 2155 335 2425
rect 355 2155 370 2425
rect 320 2140 370 2155
rect -680 1850 -630 1865
rect -680 1280 -665 1850
rect -645 1280 -630 1850
rect -680 1265 -630 1280
rect -580 1850 -530 1865
rect -580 1280 -565 1850
rect -545 1280 -530 1850
rect -580 1265 -530 1280
rect -480 1850 -430 1865
rect -480 1280 -465 1850
rect -445 1280 -430 1850
rect -480 1265 -430 1280
rect -380 1850 -330 1865
rect -380 1280 -365 1850
rect -345 1280 -330 1850
rect -380 1265 -330 1280
rect -280 1850 -230 1865
rect -280 1280 -265 1850
rect -245 1280 -230 1850
rect -280 1265 -230 1280
rect -180 1850 -130 1865
rect -180 1280 -165 1850
rect -145 1280 -130 1850
rect -180 1265 -130 1280
rect -80 1850 -30 1865
rect -80 1280 -65 1850
rect -45 1280 -30 1850
rect -80 1265 -30 1280
rect 20 1850 70 1865
rect 20 1280 35 1850
rect 55 1280 70 1850
rect 20 1265 70 1280
rect 120 1850 170 1865
rect 120 1280 135 1850
rect 155 1280 170 1850
rect 120 1265 170 1280
rect 220 1850 270 1865
rect 220 1280 235 1850
rect 255 1280 270 1850
rect 220 1265 270 1280
rect 320 1850 370 1865
rect 320 1280 335 1850
rect 355 1280 370 1850
rect 320 1265 370 1280
<< ndiffc >>
rect -665 -445 -645 125
rect -565 -445 -545 125
rect -465 -445 -445 125
rect -365 -445 -345 125
rect -265 -445 -245 125
rect -165 -445 -145 125
rect -65 -445 -45 125
rect 35 -445 55 125
rect 135 -445 155 125
rect 235 -445 255 125
rect 335 -445 355 125
<< pdiffc >>
rect -665 2655 -645 2760
rect -565 2655 -545 2760
rect -465 2655 -445 2760
rect -365 2655 -345 2760
rect -265 2655 -245 2760
rect -165 2655 -145 2760
rect -65 2655 -45 2760
rect 35 2655 55 2760
rect 135 2655 155 2760
rect 235 2655 255 2760
rect 335 2655 355 2760
rect -665 2155 -645 2425
rect -565 2155 -545 2425
rect -465 2155 -445 2425
rect -365 2155 -345 2425
rect -265 2155 -245 2425
rect -165 2155 -145 2425
rect -65 2155 -45 2425
rect 35 2155 55 2425
rect 135 2155 155 2425
rect 235 2155 255 2425
rect 335 2155 355 2425
rect -665 1280 -645 1850
rect -565 1280 -545 1850
rect -465 1280 -445 1850
rect -365 1280 -345 1850
rect -265 1280 -245 1850
rect -165 1280 -145 1850
rect -65 1280 -45 1850
rect 35 1280 55 1850
rect 135 1280 155 1850
rect 235 1280 255 1850
rect 335 1280 355 1850
<< psubdiff >>
rect -730 125 -680 140
rect -730 -445 -715 125
rect -695 -445 -680 125
rect -730 -460 -680 -445
rect 370 125 420 140
rect 370 -445 385 125
rect 405 -445 420 125
rect 370 -460 420 -445
<< nsubdiff >>
rect -730 2760 -680 2775
rect -730 2655 -715 2760
rect -695 2655 -680 2760
rect -730 2640 -680 2655
rect 370 2760 420 2775
rect 370 2655 385 2760
rect 405 2655 420 2760
rect 370 2640 420 2655
rect -730 2425 -680 2440
rect -730 2155 -715 2425
rect -695 2155 -680 2425
rect -730 2140 -680 2155
rect 370 2425 420 2440
rect 370 2155 385 2425
rect 405 2155 420 2425
rect 370 2140 420 2155
rect -730 1850 -680 1865
rect -730 1280 -715 1850
rect -695 1280 -680 1850
rect -730 1265 -680 1280
rect 370 1850 420 1865
rect 370 1280 385 1850
rect 405 1280 420 1850
rect 370 1265 420 1280
<< psubdiffcont >>
rect -715 -445 -695 125
rect 385 -445 405 125
<< nsubdiffcont >>
rect -715 2655 -695 2760
rect 385 2655 405 2760
rect -715 2155 -695 2425
rect 385 2155 405 2425
rect -715 1280 -695 1850
rect 385 1280 405 1850
<< poly >>
rect -530 2835 -480 2850
rect -530 2810 -520 2835
rect -495 2810 -480 2835
rect -630 2775 -580 2790
rect -530 2775 -480 2810
rect -430 2775 -380 2790
rect -330 2775 -280 2790
rect -230 2775 -180 2790
rect -130 2775 -80 2790
rect -30 2775 20 2790
rect 70 2775 120 2790
rect 170 2775 220 2790
rect 270 2775 320 2790
rect -630 2625 -580 2640
rect -675 2615 -580 2625
rect -675 2595 -665 2615
rect -645 2610 -580 2615
rect -530 2625 -480 2640
rect -430 2625 -380 2640
rect -330 2625 -280 2640
rect -230 2625 -180 2640
rect -130 2625 -80 2640
rect -30 2625 20 2640
rect 70 2625 120 2640
rect 170 2625 220 2640
rect -530 2610 220 2625
rect 270 2625 320 2640
rect 270 2615 365 2625
rect 270 2610 335 2615
rect -645 2595 -635 2610
rect -675 2585 -635 2595
rect 325 2595 335 2610
rect 355 2595 365 2615
rect 325 2585 365 2595
rect 375 2550 415 2560
rect 375 2535 385 2550
rect 105 2530 385 2535
rect 405 2530 415 2550
rect 105 2520 415 2530
rect 105 2495 120 2520
rect -675 2485 -635 2495
rect -675 2465 -665 2485
rect -645 2470 -635 2485
rect -430 2480 120 2495
rect -645 2465 -580 2470
rect -675 2455 -580 2465
rect -630 2440 -580 2455
rect -530 2440 -480 2455
rect -430 2440 -380 2480
rect -330 2440 -280 2480
rect -230 2440 -180 2455
rect -130 2440 -80 2455
rect -30 2440 20 2480
rect 70 2440 120 2480
rect 325 2485 365 2495
rect 325 2470 335 2485
rect 270 2465 335 2470
rect 355 2465 365 2485
rect 270 2455 365 2465
rect 170 2440 220 2455
rect 270 2440 320 2455
rect -630 2125 -580 2140
rect -530 2100 -480 2140
rect -430 2125 -380 2140
rect -330 2125 -280 2140
rect -230 2100 -180 2140
rect -130 2100 -80 2140
rect -30 2125 20 2140
rect 70 2125 120 2140
rect 170 2100 220 2140
rect 270 2125 320 2140
rect -530 2090 325 2100
rect -530 2085 295 2090
rect 285 2070 295 2085
rect 315 2070 325 2090
rect 285 2060 325 2070
rect -375 2050 65 2060
rect -375 2030 -365 2050
rect -345 2045 35 2050
rect -345 2030 -335 2045
rect -375 2020 -335 2030
rect 25 2030 35 2045
rect 55 2030 65 2050
rect 25 2020 65 2030
rect -530 1945 220 1960
rect -675 1910 -635 1920
rect -675 1890 -665 1910
rect -645 1895 -635 1910
rect -645 1890 -580 1895
rect -675 1880 -580 1890
rect -630 1865 -580 1880
rect -530 1865 -480 1945
rect -430 1865 -380 1880
rect -330 1865 -280 1880
rect -230 1865 -180 1945
rect -130 1865 -80 1945
rect -30 1865 20 1880
rect 70 1865 120 1880
rect 170 1865 220 1945
rect 325 1910 365 1920
rect 325 1895 335 1910
rect 270 1890 335 1895
rect 355 1890 365 1910
rect 270 1880 365 1890
rect 270 1865 320 1880
rect -630 1250 -580 1265
rect -725 1210 -685 1220
rect -725 1190 -715 1210
rect -695 1195 -685 1210
rect -530 1195 -480 1265
rect -695 1190 -480 1195
rect -725 1180 -480 1190
rect -430 1225 -380 1265
rect -330 1225 -280 1265
rect -230 1250 -180 1265
rect -130 1250 -80 1265
rect -30 1225 20 1265
rect 70 1225 120 1265
rect 170 1250 220 1265
rect 270 1250 320 1265
rect -430 1215 120 1225
rect -430 1210 -165 1215
rect -430 340 -415 1210
rect -175 1195 -165 1210
rect -145 1210 120 1215
rect -145 1195 -135 1210
rect -175 1185 -135 1195
rect -575 330 -415 340
rect -575 310 -565 330
rect -545 325 -415 330
rect 105 340 120 1210
rect 105 330 265 340
rect 105 325 235 330
rect -545 310 -535 325
rect -575 300 -535 310
rect 225 310 235 325
rect 255 310 265 330
rect 225 300 265 310
rect -725 250 -685 260
rect -725 230 -715 250
rect -695 235 -685 250
rect -695 230 -415 235
rect -725 220 -415 230
rect -430 195 -415 220
rect -675 185 -635 195
rect -675 165 -665 185
rect -645 170 -635 185
rect -430 180 120 195
rect -645 165 -580 170
rect -675 155 -580 165
rect -630 140 -580 155
rect -530 140 -480 155
rect -430 140 -380 180
rect -330 140 -280 180
rect -230 140 -180 155
rect -130 140 -80 155
rect -30 140 20 180
rect 70 140 120 180
rect 325 185 365 195
rect 325 170 335 185
rect 270 165 335 170
rect 355 165 365 185
rect 270 155 365 165
rect 170 140 220 155
rect 270 140 320 155
rect -630 -475 -580 -460
rect -700 -485 -660 -475
rect -700 -505 -690 -485
rect -670 -500 -660 -485
rect -530 -500 -480 -460
rect -430 -475 -380 -460
rect -330 -475 -280 -460
rect -230 -500 -180 -460
rect -130 -500 -80 -460
rect -30 -475 20 -460
rect 70 -475 120 -460
rect 170 -500 220 -460
rect 270 -475 320 -460
rect -670 -505 220 -500
rect -700 -515 220 -505
<< polycont >>
rect -520 2810 -495 2835
rect -665 2595 -645 2615
rect 335 2595 355 2615
rect 385 2530 405 2550
rect -665 2465 -645 2485
rect 335 2465 355 2485
rect 295 2070 315 2090
rect -365 2030 -345 2050
rect 35 2030 55 2050
rect -665 1890 -645 1910
rect 335 1890 355 1910
rect -715 1190 -695 1210
rect -165 1195 -145 1215
rect -565 310 -545 330
rect 235 310 255 330
rect -715 230 -695 250
rect -665 165 -645 185
rect 335 165 355 185
rect -690 -505 -670 -485
<< locali >>
rect -530 2835 -480 2850
rect -530 2820 -520 2835
rect -730 2810 -520 2820
rect -495 2810 -480 2835
rect -730 2800 -480 2810
rect -725 2760 -635 2770
rect -725 2655 -715 2760
rect -695 2655 -665 2760
rect -645 2655 -635 2760
rect -725 2645 -635 2655
rect -575 2760 -535 2770
rect -575 2655 -565 2760
rect -545 2655 -535 2760
rect -575 2645 -535 2655
rect -475 2760 -435 2770
rect -475 2655 -465 2760
rect -445 2655 -435 2760
rect -675 2615 -635 2645
rect -675 2595 -665 2615
rect -645 2595 -635 2615
rect -675 2585 -635 2595
rect -475 2615 -435 2655
rect -375 2760 -335 2770
rect -375 2655 -365 2760
rect -345 2655 -335 2760
rect -375 2645 -335 2655
rect -275 2760 -235 2770
rect -275 2655 -265 2760
rect -245 2655 -235 2760
rect -275 2615 -235 2655
rect -175 2760 -135 2770
rect -175 2655 -165 2760
rect -145 2655 -135 2760
rect -175 2645 -135 2655
rect -75 2760 -35 2770
rect -75 2655 -65 2760
rect -45 2655 -35 2760
rect -75 2615 -35 2655
rect 25 2760 65 2770
rect 25 2655 35 2760
rect 55 2655 65 2760
rect 25 2645 65 2655
rect 125 2760 165 2770
rect 125 2655 135 2760
rect 155 2655 165 2760
rect 125 2615 165 2655
rect 225 2760 265 2770
rect 225 2655 235 2760
rect 255 2655 265 2760
rect 225 2645 265 2655
rect 325 2760 415 2770
rect 325 2655 335 2760
rect 355 2655 385 2760
rect 405 2655 415 2760
rect 325 2645 415 2655
rect -475 2595 165 2615
rect -675 2485 -635 2495
rect -675 2465 -665 2485
rect -645 2465 -635 2485
rect -675 2435 -635 2465
rect -725 2425 -635 2435
rect -725 2155 -715 2425
rect -695 2155 -665 2425
rect -645 2155 -635 2425
rect -725 2145 -635 2155
rect -575 2425 -535 2435
rect -575 2155 -565 2425
rect -545 2155 -535 2425
rect -575 2000 -535 2155
rect -475 2425 -435 2595
rect -475 2155 -465 2425
rect -445 2155 -435 2425
rect -475 2145 -435 2155
rect -375 2425 -335 2435
rect -375 2155 -365 2425
rect -345 2155 -335 2425
rect -375 2060 -335 2155
rect -275 2425 -235 2595
rect -275 2155 -265 2425
rect -245 2155 -235 2425
rect -275 2145 -235 2155
rect -175 2425 -135 2435
rect -175 2155 -165 2425
rect -145 2155 -135 2425
rect -440 2050 -335 2060
rect -440 2030 -430 2050
rect -410 2040 -365 2050
rect -410 2030 -400 2040
rect -440 2020 -400 2030
rect -375 2030 -365 2040
rect -345 2030 -335 2050
rect -375 2020 -335 2030
rect -175 2010 -135 2155
rect -75 2425 -35 2595
rect -75 2155 -65 2425
rect -45 2155 -35 2425
rect -75 2145 -35 2155
rect 25 2425 65 2435
rect 25 2155 35 2425
rect 55 2155 65 2425
rect 25 2050 65 2155
rect 125 2425 165 2595
rect 325 2615 365 2645
rect 325 2595 335 2615
rect 355 2595 365 2615
rect 325 2585 365 2595
rect 375 2550 415 2560
rect 375 2530 385 2550
rect 405 2540 415 2550
rect 405 2530 420 2540
rect 375 2520 420 2530
rect 325 2485 365 2495
rect 325 2465 335 2485
rect 355 2465 365 2485
rect 325 2435 365 2465
rect 125 2155 135 2425
rect 155 2155 165 2425
rect 125 2145 165 2155
rect 225 2425 265 2435
rect 225 2155 235 2425
rect 255 2155 265 2425
rect 25 2030 35 2050
rect 55 2030 65 2050
rect 25 2020 65 2030
rect -175 2000 -165 2010
rect -575 1990 -165 2000
rect -145 2000 -135 2010
rect 225 2000 265 2155
rect 325 2425 415 2435
rect 325 2155 335 2425
rect 355 2155 385 2425
rect 405 2155 415 2425
rect 325 2145 415 2155
rect 285 2090 420 2100
rect 285 2070 295 2090
rect 315 2080 420 2090
rect 315 2070 325 2080
rect 285 2060 325 2070
rect -145 1990 265 2000
rect -575 1980 265 1990
rect -475 1920 165 1940
rect -675 1910 -635 1920
rect -675 1890 -665 1910
rect -645 1890 -635 1910
rect -675 1860 -635 1890
rect -725 1850 -635 1860
rect -725 1280 -715 1850
rect -695 1280 -665 1850
rect -645 1280 -635 1850
rect -725 1270 -635 1280
rect -575 1850 -535 1860
rect -575 1280 -565 1850
rect -545 1280 -535 1850
rect -725 1210 -685 1220
rect -725 1200 -715 1210
rect -730 1190 -715 1200
rect -695 1190 -685 1210
rect -730 1180 -685 1190
rect -575 1165 -535 1280
rect -475 1850 -435 1920
rect -275 1880 -35 1900
rect -475 1280 -465 1850
rect -445 1280 -435 1850
rect -475 1270 -435 1280
rect -375 1850 -335 1860
rect -375 1280 -365 1850
rect -345 1280 -335 1850
rect -375 1270 -335 1280
rect -275 1850 -235 1880
rect -275 1280 -265 1850
rect -245 1280 -235 1850
rect -275 1270 -235 1280
rect -175 1850 -135 1860
rect -175 1280 -165 1850
rect -145 1280 -135 1850
rect -175 1215 -135 1280
rect -75 1850 -35 1880
rect -75 1280 -65 1850
rect -45 1280 -35 1850
rect -75 1270 -35 1280
rect 25 1850 65 1860
rect 25 1280 35 1850
rect 55 1280 65 1850
rect 25 1270 65 1280
rect 125 1850 165 1920
rect 325 1910 365 1920
rect 325 1890 335 1910
rect 355 1890 365 1910
rect 325 1865 365 1890
rect 325 1860 370 1865
rect 125 1280 135 1850
rect 155 1280 165 1850
rect 125 1270 165 1280
rect 225 1850 265 1860
rect 225 1280 235 1850
rect 255 1280 265 1850
rect -175 1195 -165 1215
rect -145 1195 -135 1215
rect -175 1185 -135 1195
rect 225 1165 265 1280
rect 325 1850 415 1860
rect 325 1280 335 1850
rect 355 1280 385 1850
rect 405 1280 415 1850
rect 325 1270 415 1280
rect -575 1145 440 1165
rect -730 1090 -705 1110
rect -725 260 -705 1090
rect -575 330 -535 340
rect -575 310 -565 330
rect -545 310 -535 330
rect -725 250 -685 260
rect -725 230 -715 250
rect -695 230 -685 250
rect -725 220 -685 230
rect -675 185 -635 195
rect -675 165 -665 185
rect -645 165 -635 185
rect -675 140 -635 165
rect -680 135 -635 140
rect -725 125 -635 135
rect -725 -445 -715 125
rect -695 -445 -665 125
rect -645 -445 -635 125
rect -725 -455 -635 -445
rect -575 125 -535 310
rect -575 -445 -565 125
rect -545 -445 -535 125
rect -575 -455 -535 -445
rect -475 290 -435 300
rect -475 270 -465 290
rect -445 270 -435 290
rect -475 125 -435 270
rect -475 -445 -465 125
rect -445 -445 -435 125
rect -700 -485 -660 -475
rect -730 -505 -690 -485
rect -670 -505 -660 -485
rect -700 -515 -660 -505
rect -475 -515 -435 -445
rect -375 125 -335 135
rect -375 -445 -365 125
rect -345 -445 -335 125
rect -375 -455 -335 -445
rect -275 125 -235 135
rect -275 -445 -265 125
rect -245 -445 -235 125
rect -275 -475 -235 -445
rect -175 125 -135 1145
rect 225 330 265 340
rect 225 310 235 330
rect 255 310 265 330
rect -175 -445 -165 125
rect -145 -445 -135 125
rect -175 -455 -135 -445
rect -75 250 -35 260
rect -75 230 -65 250
rect -45 230 -35 250
rect -75 125 -35 230
rect -75 -445 -65 125
rect -45 -445 -35 125
rect -75 -475 -35 -445
rect 25 125 65 135
rect 25 -445 35 125
rect 55 -445 65 125
rect 25 -455 65 -445
rect 125 125 165 135
rect 125 -445 135 125
rect 155 -445 165 125
rect -275 -495 -35 -475
rect 125 -515 165 -445
rect 225 125 265 310
rect 225 -445 235 125
rect 255 -445 265 125
rect 225 -455 265 -445
rect 325 185 365 195
rect 325 165 335 185
rect 355 165 365 185
rect 325 135 365 165
rect 325 125 415 135
rect 325 -445 335 125
rect 355 -445 385 125
rect 405 -445 415 125
rect 325 -455 415 -445
rect -475 -535 165 -515
<< viali >>
rect -715 2655 -695 2760
rect -665 2655 -645 2760
rect -565 2655 -545 2760
rect -365 2655 -345 2760
rect -165 2655 -145 2760
rect 35 2655 55 2760
rect 235 2655 255 2760
rect 335 2655 355 2760
rect 385 2655 405 2760
rect -430 2030 -410 2050
rect -165 1990 -145 2010
rect -715 1280 -695 1850
rect -665 1280 -645 1850
rect -365 1280 -345 1850
rect 35 1280 55 1850
rect 335 1280 355 1850
rect 385 1280 405 1850
rect -715 -445 -695 125
rect -665 -445 -645 125
rect -465 270 -445 290
rect -365 -445 -345 125
rect -65 230 -45 250
rect 35 -445 55 125
rect 335 -445 355 125
rect 385 -445 405 125
<< metal1 >>
rect -730 2760 420 2770
rect -730 2655 -715 2760
rect -695 2655 -665 2760
rect -645 2655 -565 2760
rect -545 2655 -365 2760
rect -345 2655 -165 2760
rect -145 2655 35 2760
rect 55 2655 235 2760
rect 255 2655 335 2760
rect 355 2655 385 2760
rect 405 2655 420 2760
rect -730 2145 420 2655
rect -730 1860 -635 2145
rect -440 2050 -400 2060
rect -440 2030 -430 2050
rect -410 2030 -400 2050
rect -440 1930 -400 2030
rect -175 2010 -135 2020
rect -175 1990 -165 2010
rect -145 1990 -135 2010
rect -175 1930 -135 1990
rect -440 1890 -235 1930
rect -175 1890 -35 1930
rect -730 1850 -335 1860
rect -730 1280 -715 1850
rect -695 1280 -665 1850
rect -645 1280 -365 1850
rect -345 1280 -335 1850
rect -730 1270 -335 1280
rect -275 300 -235 1890
rect -475 290 -235 300
rect -475 270 -465 290
rect -445 270 -235 290
rect -475 260 -235 270
rect -75 250 -35 1890
rect 325 1860 420 2145
rect 25 1850 420 1860
rect 25 1280 35 1850
rect 55 1280 335 1850
rect 355 1280 385 1850
rect 405 1280 420 1850
rect 25 1270 420 1280
rect -75 230 -65 250
rect -45 230 -35 250
rect -75 220 -35 230
rect -725 125 415 135
rect -725 -445 -715 125
rect -695 -445 -665 125
rect -645 -445 -365 125
rect -345 -445 35 125
rect 55 -445 335 125
rect 355 -445 385 125
rect 405 -445 415 125
rect -725 -455 415 -445
<< end >>
