* SPICE3 file created from /home/madvlsi/Desktop/madvlsi/MP2/layout/csrl.ext - technology: sky130A

.subckt home/madvlsi/Desktop/madvlsi/MP2/layout/csrl VP Dn D VN CLK Q Qn
X0 VP a_80_850# a_80_1350# VP sky130_fd_pr__pfet_01v8 ad=9.5e+11p pd=5.8e+06u as=4.75e+11p ps=2.9e+06u w=950000u l=150000u
X1 Q CLK a_80_1350# VN sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X2 a_340_2000# CLK VP VP sky130_fd_pr__pfet_01v8 ad=2.375e+11p pd=2.4e+06u as=0p ps=0u w=950000u l=150000u
X3 a_340_1350# CLK VP VP sky130_fd_pr__pfet_01v8 ad=2.375e+11p pd=2.4e+06u as=0p ps=0u w=950000u l=150000u
X4 a_80_850# a_80_1350# a_80_340# VN sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=2.5e+11p ps=2.5e+06u w=1e+06u l=150000u
X5 a_80_340# CLK VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2e+12p ps=1.2e+07u w=1e+06u l=150000u
X6 a_80_1040# CLK VN VN sky130_fd_pr__nfet_01v8 ad=2.5e+11p pd=2.5e+06u as=0p ps=0u w=1e+06u l=150000u
X7 Qn CLK a_80_850# VN sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X8 a_80_850# CLK Dn VP sky130_fd_pr__pfet_01v8 ad=4.75e+11p pd=2.9e+06u as=4.75e+11p ps=2.9e+06u w=950000u l=150000u
X9 a_80_1350# a_80_850# a_80_1040# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VN Qn Q VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_80_1350# CLK D VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.75e+11p ps=2.9e+06u w=950000u l=150000u
X12 VN Q Qn VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Qn Q a_340_2000# VP sky130_fd_pr__pfet_01v8 ad=4.75e+11p pd=2.9e+06u as=0p ps=0u w=950000u l=150000u
X14 VP a_80_1350# a_80_850# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=950000u l=150000u
X15 Q Qn a_340_1350# VP sky130_fd_pr__pfet_01v8 ad=4.75e+11p pd=2.9e+06u as=0p ps=0u w=950000u l=150000u
.ends

