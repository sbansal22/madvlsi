magic
tech sky130A
timestamp 1615761100
<< nwell >>
rect -70 2430 1320 4320
<< nmos >>
rect 50 1000 100 1600
rect 150 1000 200 1600
rect 250 1000 300 1600
rect 350 1000 400 1600
rect 550 1000 600 1600
rect 650 1000 700 1600
rect 850 1000 900 1600
rect 950 1000 1000 1600
rect 1050 1000 1100 1600
rect 1150 1000 1200 1600
rect 50 -300 100 300
rect 150 -300 200 300
rect 250 -300 300 300
rect 350 -300 400 300
rect 550 -300 600 300
rect 650 -300 700 300
rect 850 -300 900 300
rect 950 -300 1000 300
rect 1050 -300 1100 300
rect 1150 -300 1200 300
<< pmos >>
rect 50 3700 100 4300
rect 150 3700 200 4300
rect 250 3700 300 4300
rect 450 3700 500 4300
rect 550 3700 600 4300
rect 650 3700 700 4300
rect 750 3700 800 4300
rect 950 3700 1000 4300
rect 1050 3700 1100 4300
rect 1150 3700 1200 4300
rect 50 2450 100 3050
rect 150 2450 200 3050
rect 250 2450 300 3050
rect 350 2450 400 3050
rect 550 2450 600 3050
rect 650 2450 700 3050
rect 850 2450 900 3050
rect 950 2450 1000 3050
rect 1050 2450 1100 3050
rect 1150 2450 1200 3050
<< ndiff >>
rect 0 1585 50 1600
rect 0 1015 15 1585
rect 35 1015 50 1585
rect 0 1000 50 1015
rect 100 1585 150 1600
rect 100 1015 115 1585
rect 135 1015 150 1585
rect 100 1000 150 1015
rect 200 1585 250 1600
rect 200 1015 215 1585
rect 235 1015 250 1585
rect 200 1000 250 1015
rect 300 1585 350 1600
rect 300 1015 315 1585
rect 335 1015 350 1585
rect 300 1000 350 1015
rect 400 1585 450 1600
rect 400 1015 415 1585
rect 435 1015 450 1585
rect 400 1000 450 1015
rect 500 1585 550 1600
rect 500 1015 515 1585
rect 535 1015 550 1585
rect 500 1000 550 1015
rect 600 1585 650 1600
rect 600 1015 615 1585
rect 635 1015 650 1585
rect 600 1000 650 1015
rect 700 1585 750 1600
rect 700 1015 715 1585
rect 735 1015 750 1585
rect 700 1000 750 1015
rect 800 1585 850 1600
rect 800 1015 815 1585
rect 835 1015 850 1585
rect 800 1000 850 1015
rect 900 1585 950 1600
rect 900 1015 915 1585
rect 935 1015 950 1585
rect 900 1000 950 1015
rect 1000 1585 1050 1600
rect 1000 1015 1015 1585
rect 1035 1015 1050 1585
rect 1000 1000 1050 1015
rect 1100 1585 1150 1600
rect 1100 1015 1115 1585
rect 1135 1015 1150 1585
rect 1100 1000 1150 1015
rect 1200 1585 1250 1600
rect 1200 1015 1215 1585
rect 1235 1015 1250 1585
rect 1200 1000 1250 1015
rect 0 285 50 300
rect 0 -285 15 285
rect 35 -285 50 285
rect 0 -300 50 -285
rect 100 285 150 300
rect 100 -285 115 285
rect 135 -285 150 285
rect 100 -300 150 -285
rect 200 285 250 300
rect 200 -285 215 285
rect 235 -285 250 285
rect 200 -300 250 -285
rect 300 285 350 300
rect 300 -285 315 285
rect 335 -285 350 285
rect 300 -300 350 -285
rect 400 285 450 300
rect 400 -285 415 285
rect 435 -285 450 285
rect 400 -300 450 -285
rect 500 285 550 300
rect 500 -285 515 285
rect 535 -285 550 285
rect 500 -300 550 -285
rect 600 285 650 300
rect 600 -285 615 285
rect 635 -285 650 285
rect 600 -300 650 -285
rect 700 285 750 300
rect 700 -285 715 285
rect 735 -285 750 285
rect 700 -300 750 -285
rect 800 285 850 300
rect 800 -285 815 285
rect 835 -285 850 285
rect 800 -300 850 -285
rect 900 285 950 300
rect 900 -285 915 285
rect 935 -285 950 285
rect 900 -300 950 -285
rect 1000 285 1050 300
rect 1000 -285 1015 285
rect 1035 -285 1050 285
rect 1000 -300 1050 -285
rect 1100 285 1150 300
rect 1100 -285 1115 285
rect 1135 -285 1150 285
rect 1100 -300 1150 -285
rect 1200 285 1250 300
rect 1200 -285 1215 285
rect 1235 -285 1250 285
rect 1200 -300 1250 -285
<< pdiff >>
rect 0 4285 50 4300
rect 0 3715 15 4285
rect 35 3715 50 4285
rect 0 3700 50 3715
rect 100 4285 150 4300
rect 100 3715 115 4285
rect 135 3715 150 4285
rect 100 3700 150 3715
rect 200 4285 250 4300
rect 200 3715 215 4285
rect 235 3715 250 4285
rect 200 3700 250 3715
rect 300 4285 350 4300
rect 300 3715 315 4285
rect 335 3715 350 4285
rect 300 3700 350 3715
rect 400 4285 450 4300
rect 400 3715 415 4285
rect 435 3715 450 4285
rect 400 3700 450 3715
rect 500 4285 550 4300
rect 500 3715 515 4285
rect 535 3715 550 4285
rect 500 3700 550 3715
rect 600 4285 650 4300
rect 600 3715 615 4285
rect 635 3715 650 4285
rect 600 3700 650 3715
rect 700 4285 750 4300
rect 700 3715 715 4285
rect 735 3715 750 4285
rect 700 3700 750 3715
rect 800 4285 850 4300
rect 800 3715 815 4285
rect 835 3715 850 4285
rect 800 3700 850 3715
rect 900 4285 950 4300
rect 900 3715 915 4285
rect 935 3715 950 4285
rect 900 3700 950 3715
rect 1000 4285 1050 4300
rect 1000 3715 1015 4285
rect 1035 3715 1050 4285
rect 1000 3700 1050 3715
rect 1100 4285 1150 4300
rect 1100 3715 1115 4285
rect 1135 3715 1150 4285
rect 1100 3700 1150 3715
rect 1200 4285 1250 4300
rect 1200 3715 1215 4285
rect 1235 3715 1250 4285
rect 1200 3700 1250 3715
rect 0 3035 50 3050
rect 0 2465 15 3035
rect 35 2465 50 3035
rect 0 2450 50 2465
rect 100 3035 150 3050
rect 100 2465 115 3035
rect 135 2465 150 3035
rect 100 2450 150 2465
rect 200 3035 250 3050
rect 200 2465 215 3035
rect 235 2465 250 3035
rect 200 2450 250 2465
rect 300 3035 350 3050
rect 300 2465 315 3035
rect 335 2465 350 3035
rect 300 2450 350 2465
rect 400 3035 450 3050
rect 400 2465 415 3035
rect 435 2465 450 3035
rect 400 2450 450 2465
rect 500 3035 550 3050
rect 500 2465 515 3035
rect 535 2465 550 3035
rect 500 2450 550 2465
rect 600 3035 650 3050
rect 600 2465 615 3035
rect 635 2465 650 3035
rect 600 2450 650 2465
rect 700 3035 750 3050
rect 700 2465 715 3035
rect 735 2465 750 3035
rect 700 2450 750 2465
rect 800 3035 850 3050
rect 800 2465 815 3035
rect 835 2465 850 3035
rect 800 2450 850 2465
rect 900 3035 950 3050
rect 900 2465 915 3035
rect 935 2465 950 3035
rect 900 2450 950 2465
rect 1000 3035 1050 3050
rect 1000 2465 1015 3035
rect 1035 2465 1050 3035
rect 1000 2450 1050 2465
rect 1100 3035 1150 3050
rect 1100 2465 1115 3035
rect 1135 2465 1150 3035
rect 1100 2450 1150 2465
rect 1200 3035 1250 3050
rect 1200 2465 1215 3035
rect 1235 2465 1250 3035
rect 1200 2450 1250 2465
<< ndiffc >>
rect 15 1015 35 1585
rect 115 1015 135 1585
rect 215 1015 235 1585
rect 315 1015 335 1585
rect 415 1015 435 1585
rect 515 1015 535 1585
rect 615 1015 635 1585
rect 715 1015 735 1585
rect 815 1015 835 1585
rect 915 1015 935 1585
rect 1015 1015 1035 1585
rect 1115 1015 1135 1585
rect 1215 1015 1235 1585
rect 15 -285 35 285
rect 115 -285 135 285
rect 215 -285 235 285
rect 315 -285 335 285
rect 415 -285 435 285
rect 515 -285 535 285
rect 615 -285 635 285
rect 715 -285 735 285
rect 815 -285 835 285
rect 915 -285 935 285
rect 1015 -285 1035 285
rect 1115 -285 1135 285
rect 1215 -285 1235 285
<< pdiffc >>
rect 15 3715 35 4285
rect 115 3715 135 4285
rect 215 3715 235 4285
rect 315 3715 335 4285
rect 415 3715 435 4285
rect 515 3715 535 4285
rect 615 3715 635 4285
rect 715 3715 735 4285
rect 815 3715 835 4285
rect 915 3715 935 4285
rect 1015 3715 1035 4285
rect 1115 3715 1135 4285
rect 1215 3715 1235 4285
rect 15 2465 35 3035
rect 115 2465 135 3035
rect 215 2465 235 3035
rect 315 2465 335 3035
rect 415 2465 435 3035
rect 515 2465 535 3035
rect 615 2465 635 3035
rect 715 2465 735 3035
rect 815 2465 835 3035
rect 915 2465 935 3035
rect 1015 2465 1035 3035
rect 1115 2465 1135 3035
rect 1215 2465 1235 3035
<< psubdiff >>
rect -50 1585 0 1600
rect -50 1015 -35 1585
rect -15 1015 0 1585
rect -50 1000 0 1015
rect 1250 1585 1300 1600
rect 1250 1015 1265 1585
rect 1285 1015 1300 1585
rect 1250 1000 1300 1015
rect -50 285 0 300
rect -50 -285 -35 285
rect -15 -285 0 285
rect -50 -300 0 -285
rect 1250 285 1300 300
rect 1250 -285 1265 285
rect 1285 -285 1300 285
rect 1250 -300 1300 -285
<< nsubdiff >>
rect -50 4285 0 4300
rect -50 3715 -35 4285
rect -15 3715 0 4285
rect -50 3700 0 3715
rect 1250 4285 1300 4300
rect 1250 3715 1265 4285
rect 1285 3715 1300 4285
rect 1250 3700 1300 3715
rect -50 3035 0 3050
rect -50 2465 -35 3035
rect -15 2465 0 3035
rect -50 2450 0 2465
rect 1250 3035 1300 3050
rect 1250 2465 1265 3035
rect 1285 2465 1300 3035
rect 1250 2450 1300 2465
<< psubdiffcont >>
rect -35 1015 -15 1585
rect 1265 1015 1285 1585
rect -35 -285 -15 285
rect 1265 -285 1285 285
<< nsubdiffcont >>
rect -35 3715 -15 4285
rect 1265 3715 1285 4285
rect -35 2465 -15 3035
rect 1265 2465 1285 3035
<< poly >>
rect 50 4300 100 4315
rect 150 4300 200 4315
rect 250 4300 300 4315
rect 450 4300 500 4315
rect 550 4300 600 4315
rect 650 4300 700 4315
rect 750 4300 800 4315
rect 950 4300 1000 4315
rect 1050 4300 1100 4315
rect 1150 4300 1200 4315
rect 50 3685 100 3700
rect 5 3675 100 3685
rect 5 3655 15 3675
rect 35 3670 100 3675
rect 150 3685 200 3700
rect 250 3685 300 3700
rect 450 3685 500 3700
rect 550 3685 600 3700
rect 650 3685 700 3700
rect 750 3685 800 3700
rect 950 3685 1000 3700
rect 1050 3685 1100 3700
rect 150 3670 1100 3685
rect 1150 3685 1200 3700
rect 1150 3675 1245 3685
rect 1150 3670 1215 3675
rect 35 3655 45 3670
rect 5 3645 45 3655
rect 150 3645 165 3670
rect 70 3635 165 3645
rect 70 3615 80 3635
rect 100 3630 165 3635
rect 1085 3645 1100 3670
rect 1205 3655 1215 3670
rect 1235 3655 1245 3675
rect 1205 3645 1245 3655
rect 1085 3635 1180 3645
rect 1085 3630 1150 3635
rect 100 3615 110 3630
rect 70 3605 110 3615
rect 1140 3615 1150 3630
rect 1170 3615 1180 3635
rect 1140 3605 1180 3615
rect 405 3120 845 3130
rect 405 3105 415 3120
rect 105 3095 145 3105
rect 105 3080 115 3095
rect 50 3075 115 3080
rect 135 3080 145 3095
rect 385 3100 415 3105
rect 435 3115 815 3120
rect 435 3100 445 3115
rect 385 3090 445 3100
rect 805 3100 815 3115
rect 835 3105 845 3120
rect 835 3100 865 3105
rect 805 3090 865 3100
rect 385 3080 400 3090
rect 850 3080 865 3090
rect 1105 3095 1145 3105
rect 1105 3080 1115 3095
rect 135 3075 200 3080
rect 50 3065 200 3075
rect 50 3050 100 3065
rect 150 3050 200 3065
rect 250 3065 400 3080
rect 250 3050 300 3065
rect 350 3050 400 3065
rect 550 3065 700 3080
rect 550 3050 600 3065
rect 650 3050 700 3065
rect 850 3065 1000 3080
rect 850 3050 900 3065
rect 950 3050 1000 3065
rect 1050 3075 1115 3080
rect 1135 3080 1145 3095
rect 1135 3075 1200 3080
rect 1050 3065 1200 3075
rect 1050 3050 1100 3065
rect 1150 3050 1200 3065
rect 50 2435 100 2450
rect 150 2435 200 2450
rect 250 1735 300 2450
rect 350 2435 400 2450
rect 550 1775 600 2450
rect 650 2435 700 2450
rect 850 2435 900 2450
rect 950 2435 1000 2450
rect 1050 2435 1100 2450
rect 1150 2435 1200 2450
rect 550 1755 565 1775
rect 585 1755 600 1775
rect 550 1745 600 1755
rect 250 1715 265 1735
rect 285 1720 300 1735
rect 925 1735 965 1745
rect 925 1720 935 1735
rect 285 1715 935 1720
rect 955 1715 965 1735
rect 250 1705 965 1715
rect 985 1685 1210 1695
rect 985 1680 1180 1685
rect 405 1670 445 1680
rect 405 1655 415 1670
rect 105 1645 145 1655
rect 105 1630 115 1645
rect 50 1625 115 1630
rect 135 1630 145 1645
rect 385 1650 415 1655
rect 435 1655 445 1670
rect 805 1670 845 1680
rect 805 1655 815 1670
rect 435 1650 815 1655
rect 835 1655 845 1670
rect 835 1650 865 1655
rect 385 1640 865 1650
rect 385 1630 400 1640
rect 135 1625 200 1630
rect 50 1615 200 1625
rect 50 1600 100 1615
rect 150 1600 200 1615
rect 250 1615 400 1630
rect 250 1600 300 1615
rect 350 1600 400 1615
rect 550 1600 600 1640
rect 650 1600 700 1640
rect 850 1630 865 1640
rect 985 1630 1000 1680
rect 1170 1665 1180 1680
rect 1200 1665 1210 1685
rect 1170 1655 1210 1665
rect 1105 1645 1145 1655
rect 1105 1630 1115 1645
rect 850 1615 1000 1630
rect 850 1600 900 1615
rect 950 1600 1000 1615
rect 1050 1625 1115 1630
rect 1135 1630 1145 1645
rect 1135 1625 1200 1630
rect 1050 1615 1200 1625
rect 1050 1600 1100 1615
rect 1150 1600 1200 1615
rect 50 985 100 1000
rect 150 985 200 1000
rect 250 985 300 1000
rect 350 985 400 1000
rect 550 985 600 1000
rect 650 985 700 1000
rect 850 985 900 1000
rect 950 985 1000 1000
rect 1050 985 1100 1000
rect 1150 985 1200 1000
rect 550 970 700 985
rect 405 370 445 380
rect 405 355 415 370
rect 105 345 145 355
rect 105 330 115 345
rect 50 325 115 330
rect 135 330 145 345
rect 385 350 415 355
rect 435 355 445 370
rect 805 370 845 380
rect 805 355 815 370
rect 435 350 815 355
rect 835 355 845 370
rect 835 350 865 355
rect 385 340 865 350
rect 385 330 400 340
rect 135 325 200 330
rect 50 315 200 325
rect 50 300 100 315
rect 150 300 200 315
rect 250 315 400 330
rect 850 330 865 340
rect 1105 345 1145 355
rect 1105 330 1115 345
rect 850 315 1000 330
rect 250 300 300 315
rect 350 300 400 315
rect 550 300 600 315
rect 650 300 700 315
rect 850 300 900 315
rect 950 300 1000 315
rect 1050 325 1115 330
rect 1135 330 1145 345
rect 1135 325 1200 330
rect 1050 315 1200 325
rect 1050 300 1100 315
rect 1150 300 1200 315
rect 50 -315 100 -300
rect 150 -315 200 -300
rect 250 -315 300 -300
rect 350 -315 400 -300
rect 550 -315 600 -300
rect 650 -315 700 -300
rect 850 -315 900 -300
rect 950 -315 1000 -300
rect 1050 -315 1100 -300
rect 1150 -315 1200 -300
rect 550 -325 700 -315
rect 550 -330 615 -325
rect 605 -345 615 -330
rect 635 -330 700 -325
rect 635 -345 645 -330
rect 605 -355 645 -345
<< polycont >>
rect 15 3655 35 3675
rect 80 3615 100 3635
rect 1215 3655 1235 3675
rect 1150 3615 1170 3635
rect 115 3075 135 3095
rect 415 3100 435 3120
rect 815 3100 835 3120
rect 1115 3075 1135 3095
rect 565 1755 585 1775
rect 265 1715 285 1735
rect 935 1715 955 1735
rect 115 1625 135 1645
rect 415 1650 435 1670
rect 815 1650 835 1670
rect 1180 1665 1200 1685
rect 1115 1625 1135 1645
rect 115 325 135 345
rect 415 350 435 370
rect 815 350 835 370
rect 1115 325 1135 345
rect 615 -345 635 -325
<< locali >>
rect -45 4285 45 4295
rect -45 3715 -35 4285
rect -15 3715 15 4285
rect 35 3715 45 4285
rect -45 3705 45 3715
rect 5 3675 45 3705
rect 5 3655 15 3675
rect 35 3655 45 3675
rect 5 3645 45 3655
rect 105 4285 145 4295
rect 105 3715 115 4285
rect 135 3715 145 4285
rect 105 3645 145 3715
rect 205 4285 245 4295
rect 205 3715 215 4285
rect 235 3715 245 4285
rect 205 3700 245 3715
rect 305 4285 345 4295
rect 305 3715 315 4285
rect 335 3715 345 4285
rect 70 3635 145 3645
rect 70 3625 80 3635
rect -70 3615 80 3625
rect 100 3615 145 3635
rect -70 3605 145 3615
rect 305 3510 345 3715
rect 405 4285 445 4295
rect 405 3715 415 4285
rect 435 3715 445 4285
rect 405 3565 445 3715
rect 505 4285 545 4295
rect 505 3715 515 4285
rect 535 3715 545 4285
rect 505 3705 545 3715
rect 605 4285 645 4295
rect 605 3715 615 4285
rect 635 3715 645 4285
rect 605 3605 645 3715
rect 705 4285 745 4295
rect 705 3715 715 4285
rect 735 3715 745 4285
rect 705 3705 745 3715
rect 805 4285 845 4295
rect 805 3715 815 4285
rect 835 3715 845 4285
rect 805 3565 845 3715
rect 405 3545 845 3565
rect 905 4285 945 4295
rect 905 3715 915 4285
rect 935 3715 945 4285
rect 905 3510 945 3715
rect 1005 4285 1045 4295
rect 1005 3715 1015 4285
rect 1035 3715 1045 4285
rect 1005 3705 1045 3715
rect 1105 4285 1145 4295
rect 1105 3715 1115 4285
rect 1135 3715 1145 4285
rect 1105 3645 1145 3715
rect 1205 4285 1295 4295
rect 1205 3715 1215 4285
rect 1235 3715 1265 4285
rect 1285 3715 1295 4285
rect 1205 3705 1295 3715
rect 1205 3675 1245 3705
rect 1205 3655 1215 3675
rect 1235 3655 1245 3675
rect 1205 3645 1245 3655
rect 1105 3635 1180 3645
rect 1105 3615 1150 3635
rect 1170 3615 1180 3635
rect 1105 3605 1180 3615
rect 305 3490 945 3510
rect 405 3120 445 3130
rect 105 3095 145 3105
rect 105 3085 115 3095
rect 5 3075 115 3085
rect 135 3075 145 3095
rect 5 3065 145 3075
rect 405 3100 415 3120
rect 435 3100 445 3120
rect 5 3045 45 3065
rect -45 3035 45 3045
rect -45 2465 -35 3035
rect -15 2465 15 3035
rect 35 2465 45 3035
rect -45 2455 45 2465
rect 105 3035 145 3045
rect 105 2465 115 3035
rect 135 2465 145 3035
rect 105 2455 145 2465
rect 205 3035 245 3045
rect 205 2465 215 3035
rect 235 2465 245 3035
rect 205 2455 245 2465
rect 305 3035 345 3045
rect 305 2465 315 3035
rect 335 2465 345 3035
rect 305 2430 345 2465
rect 405 3035 445 3100
rect 805 3120 845 3130
rect 805 3100 815 3120
rect 835 3100 845 3120
rect 405 2465 415 3035
rect 435 2465 445 3035
rect 405 2455 445 2465
rect 505 3035 545 3045
rect 505 2465 515 3035
rect 535 2465 545 3035
rect 505 2430 545 2465
rect 605 3035 645 3045
rect 605 2465 615 3035
rect 635 2465 645 3035
rect 605 2455 645 2465
rect 705 3035 745 3045
rect 705 2465 715 3035
rect 735 2465 745 3035
rect 705 2430 745 2465
rect 805 3035 845 3100
rect 1105 3095 1145 3105
rect 1105 3075 1115 3095
rect 1135 3085 1145 3095
rect 1135 3075 1245 3085
rect 1105 3065 1245 3075
rect 1205 3045 1245 3065
rect 805 2465 815 3035
rect 835 2465 845 3035
rect 805 2455 845 2465
rect 905 3035 945 3045
rect 905 2465 915 3035
rect 935 2465 945 3035
rect 905 2430 945 2465
rect 1005 3035 1045 3045
rect 1005 2465 1015 3035
rect 1035 2465 1045 3035
rect 1005 2455 1045 2465
rect 1105 3035 1145 3045
rect 1105 2465 1115 3035
rect 1135 2465 1145 3035
rect 1105 2455 1145 2465
rect 1205 3035 1295 3045
rect 1205 2465 1215 3035
rect 1235 2465 1265 3035
rect 1285 2465 1295 3035
rect 1205 2455 1295 2465
rect 305 2410 945 2430
rect 550 1775 1300 1785
rect 550 1755 565 1775
rect 585 1765 1300 1775
rect 585 1755 645 1765
rect 550 1745 645 1755
rect 250 1735 300 1745
rect 250 1725 265 1735
rect 205 1715 265 1725
rect 285 1715 300 1735
rect 205 1705 300 1715
rect 105 1645 145 1655
rect 105 1635 115 1645
rect 5 1625 115 1635
rect 135 1625 145 1645
rect 5 1615 145 1625
rect 5 1595 45 1615
rect -45 1585 45 1595
rect -45 1015 -35 1585
rect -15 1015 15 1585
rect 35 1015 45 1585
rect -45 1005 45 1015
rect 105 1585 145 1595
rect 105 1015 115 1585
rect 135 1015 145 1585
rect 105 1005 145 1015
rect 205 1585 245 1705
rect 405 1670 445 1680
rect 405 1650 415 1670
rect 435 1650 445 1670
rect 205 1015 215 1585
rect 235 1015 245 1585
rect 205 1005 245 1015
rect 305 1585 345 1595
rect 305 1015 315 1585
rect 335 1015 345 1585
rect 305 1005 345 1015
rect 405 1585 445 1650
rect 405 1015 415 1585
rect 435 1015 445 1585
rect 405 1005 445 1015
rect 505 1585 545 1595
rect 505 1015 515 1585
rect 535 1015 545 1585
rect 505 1005 545 1015
rect 605 1585 645 1745
rect 925 1735 965 1745
rect 925 1715 935 1735
rect 955 1725 965 1735
rect 955 1715 1045 1725
rect 925 1705 1045 1715
rect 805 1670 845 1680
rect 805 1650 815 1670
rect 835 1650 845 1670
rect 605 1015 615 1585
rect 635 1015 645 1585
rect 605 1005 645 1015
rect 705 1585 745 1595
rect 705 1015 715 1585
rect 735 1015 745 1585
rect 705 1005 745 1015
rect 805 1585 845 1650
rect 805 1015 815 1585
rect 835 1015 845 1585
rect 805 1005 845 1015
rect 905 1585 945 1595
rect 905 1015 915 1585
rect 935 1015 945 1585
rect 905 1005 945 1015
rect 1005 1585 1045 1705
rect 1170 1685 1300 1695
rect 1170 1665 1180 1685
rect 1200 1675 1300 1685
rect 1200 1665 1210 1675
rect 1170 1655 1210 1665
rect 1105 1645 1145 1655
rect 1105 1625 1115 1645
rect 1135 1635 1145 1645
rect 1135 1625 1245 1635
rect 1105 1615 1245 1625
rect 1205 1595 1245 1615
rect 1005 1015 1015 1585
rect 1035 1015 1045 1585
rect 1005 1005 1045 1015
rect 1105 1585 1145 1595
rect 1105 1015 1115 1585
rect 1135 1015 1145 1585
rect 1105 1005 1145 1015
rect 1205 1585 1295 1595
rect 1205 1015 1215 1585
rect 1235 1015 1265 1585
rect 1285 1015 1295 1585
rect 1205 1005 1295 1015
rect 305 575 945 595
rect 105 345 145 355
rect 105 335 115 345
rect 5 325 115 335
rect 135 325 145 345
rect 5 315 145 325
rect 5 295 45 315
rect -45 285 45 295
rect -45 -285 -35 285
rect -15 -285 15 285
rect 35 -285 45 285
rect -45 -295 45 -285
rect 105 285 145 295
rect 105 -285 115 285
rect 135 -285 145 285
rect 105 -295 145 -285
rect 205 285 245 295
rect 205 -285 215 285
rect 235 -285 245 285
rect 205 -295 245 -285
rect 305 285 345 575
rect 305 -285 315 285
rect 335 -285 345 285
rect 305 -295 345 -285
rect 405 370 445 380
rect 405 350 415 370
rect 435 350 445 370
rect 405 285 445 350
rect 405 -285 415 285
rect 435 -285 445 285
rect 405 -295 445 -285
rect 505 285 545 575
rect 505 -285 515 285
rect 535 -285 545 285
rect 505 -295 545 -285
rect 605 285 645 475
rect 605 -285 615 285
rect 635 -285 645 285
rect 605 -295 645 -285
rect 705 285 745 575
rect 705 -285 715 285
rect 735 -285 745 285
rect 705 -295 745 -285
rect 805 370 845 380
rect 805 350 815 370
rect 835 350 845 370
rect 805 285 845 350
rect 805 -285 815 285
rect 835 -285 845 285
rect 805 -295 845 -285
rect 905 285 945 575
rect 1105 345 1145 355
rect 1105 325 1115 345
rect 1135 335 1145 345
rect 1135 325 1245 335
rect 1105 315 1245 325
rect 1205 295 1245 315
rect 905 -285 915 285
rect 935 -285 945 285
rect 905 -295 945 -285
rect 1005 285 1045 295
rect 1005 -285 1015 285
rect 1035 -285 1045 285
rect 1005 -295 1045 -285
rect 1105 285 1145 295
rect 1105 -285 1115 285
rect 1135 -285 1145 285
rect 1105 -295 1145 -285
rect 1205 285 1295 295
rect 1205 -285 1215 285
rect 1235 -285 1265 285
rect 1285 -285 1295 285
rect 1205 -295 1295 -285
rect 605 -325 645 -315
rect 605 -345 615 -325
rect 635 -345 1300 -325
rect 605 -355 645 -345
<< end >>
