magic
tech sky130A
timestamp 1615929122
<< nwell >>
rect -750 1230 440 2795
<< nmos >>
rect -630 -460 -580 140
rect -530 -460 -480 140
rect -430 -460 -380 140
rect -330 -460 -280 140
rect -230 -460 -180 140
rect -130 -460 -80 140
rect -30 -460 20 140
rect 70 -460 120 140
rect 170 -460 220 140
rect 270 -460 320 140
<< pmos >>
rect -630 2625 -580 2775
rect -530 2625 -480 2775
rect -430 2625 -380 2775
rect -330 2625 -280 2775
rect -230 2625 -180 2775
rect -130 2625 -80 2775
rect -30 2625 20 2775
rect 70 2625 120 2775
rect 170 2625 220 2775
rect 270 2625 320 2775
rect -630 2125 -580 2425
rect -530 2125 -480 2425
rect -430 2125 -380 2425
rect -330 2125 -280 2425
rect -230 2125 -180 2425
rect -130 2125 -80 2425
rect -30 2125 20 2425
rect 70 2125 120 2425
rect 170 2125 220 2425
rect 270 2125 320 2425
rect -630 1250 -580 1850
rect -530 1250 -480 1850
rect -430 1250 -380 1850
rect -330 1250 -280 1850
rect -230 1250 -180 1850
rect -130 1250 -80 1850
rect -30 1250 20 1850
rect 70 1250 120 1850
rect 170 1250 220 1850
rect 270 1250 320 1850
<< ndiff >>
rect -680 125 -630 140
rect -680 -445 -665 125
rect -645 -445 -630 125
rect -680 -460 -630 -445
rect -580 125 -530 140
rect -580 -445 -565 125
rect -545 -445 -530 125
rect -580 -460 -530 -445
rect -480 125 -430 140
rect -480 -445 -465 125
rect -445 -445 -430 125
rect -480 -460 -430 -445
rect -380 125 -330 140
rect -380 -445 -365 125
rect -345 -445 -330 125
rect -380 -460 -330 -445
rect -280 125 -230 140
rect -280 -445 -265 125
rect -245 -445 -230 125
rect -280 -460 -230 -445
rect -180 125 -130 140
rect -180 -445 -165 125
rect -145 -445 -130 125
rect -180 -460 -130 -445
rect -80 125 -30 140
rect -80 -445 -65 125
rect -45 -445 -30 125
rect -80 -460 -30 -445
rect 20 125 70 140
rect 20 -445 35 125
rect 55 -445 70 125
rect 20 -460 70 -445
rect 120 125 170 140
rect 120 -445 135 125
rect 155 -445 170 125
rect 120 -460 170 -445
rect 220 125 270 140
rect 220 -445 235 125
rect 255 -445 270 125
rect 220 -460 270 -445
rect 320 125 370 140
rect 320 -445 335 125
rect 355 -445 370 125
rect 320 -460 370 -445
<< pdiff >>
rect -680 2760 -630 2775
rect -680 2640 -665 2760
rect -645 2640 -630 2760
rect -680 2625 -630 2640
rect -580 2760 -530 2775
rect -580 2640 -565 2760
rect -545 2640 -530 2760
rect -580 2625 -530 2640
rect -480 2760 -430 2775
rect -480 2640 -465 2760
rect -445 2640 -430 2760
rect -480 2625 -430 2640
rect -380 2760 -330 2775
rect -380 2640 -365 2760
rect -345 2640 -330 2760
rect -380 2625 -330 2640
rect -280 2760 -230 2775
rect -280 2640 -265 2760
rect -245 2640 -230 2760
rect -280 2625 -230 2640
rect -180 2760 -130 2775
rect -180 2640 -165 2760
rect -145 2640 -130 2760
rect -180 2625 -130 2640
rect -80 2760 -30 2775
rect -80 2640 -65 2760
rect -45 2640 -30 2760
rect -80 2625 -30 2640
rect 20 2760 70 2775
rect 20 2640 35 2760
rect 55 2640 70 2760
rect 20 2625 70 2640
rect 120 2760 170 2775
rect 120 2640 135 2760
rect 155 2640 170 2760
rect 120 2625 170 2640
rect 220 2760 270 2775
rect 220 2640 235 2760
rect 255 2640 270 2760
rect 220 2625 270 2640
rect 320 2760 370 2775
rect 320 2640 335 2760
rect 355 2640 370 2760
rect 320 2625 370 2640
rect -680 2410 -630 2425
rect -680 2140 -665 2410
rect -645 2140 -630 2410
rect -680 2125 -630 2140
rect -580 2410 -530 2425
rect -580 2140 -565 2410
rect -545 2140 -530 2410
rect -580 2125 -530 2140
rect -480 2410 -430 2425
rect -480 2140 -465 2410
rect -445 2140 -430 2410
rect -480 2125 -430 2140
rect -380 2410 -330 2425
rect -380 2140 -365 2410
rect -345 2140 -330 2410
rect -380 2125 -330 2140
rect -280 2410 -230 2425
rect -280 2140 -265 2410
rect -245 2140 -230 2410
rect -280 2125 -230 2140
rect -180 2410 -130 2425
rect -180 2140 -165 2410
rect -145 2140 -130 2410
rect -180 2125 -130 2140
rect -80 2410 -30 2425
rect -80 2140 -65 2410
rect -45 2140 -30 2410
rect -80 2125 -30 2140
rect 20 2410 70 2425
rect 20 2140 35 2410
rect 55 2140 70 2410
rect 20 2125 70 2140
rect 120 2410 170 2425
rect 120 2140 135 2410
rect 155 2140 170 2410
rect 120 2125 170 2140
rect 220 2410 270 2425
rect 220 2140 235 2410
rect 255 2140 270 2410
rect 220 2125 270 2140
rect 320 2410 370 2425
rect 320 2140 335 2410
rect 355 2140 370 2410
rect 320 2125 370 2140
rect -680 1835 -630 1850
rect -680 1265 -665 1835
rect -645 1265 -630 1835
rect -680 1250 -630 1265
rect -580 1835 -530 1850
rect -580 1265 -565 1835
rect -545 1265 -530 1835
rect -580 1250 -530 1265
rect -480 1835 -430 1850
rect -480 1265 -465 1835
rect -445 1265 -430 1835
rect -480 1250 -430 1265
rect -380 1835 -330 1850
rect -380 1265 -365 1835
rect -345 1265 -330 1835
rect -380 1250 -330 1265
rect -280 1835 -230 1850
rect -280 1265 -265 1835
rect -245 1265 -230 1835
rect -280 1250 -230 1265
rect -180 1835 -130 1850
rect -180 1265 -165 1835
rect -145 1265 -130 1835
rect -180 1250 -130 1265
rect -80 1835 -30 1850
rect -80 1265 -65 1835
rect -45 1265 -30 1835
rect -80 1250 -30 1265
rect 20 1835 70 1850
rect 20 1265 35 1835
rect 55 1265 70 1835
rect 20 1250 70 1265
rect 120 1835 170 1850
rect 120 1265 135 1835
rect 155 1265 170 1835
rect 120 1250 170 1265
rect 220 1835 270 1850
rect 220 1265 235 1835
rect 255 1265 270 1835
rect 220 1250 270 1265
rect 320 1835 370 1850
rect 320 1265 335 1835
rect 355 1265 370 1835
rect 320 1250 370 1265
<< ndiffc >>
rect -665 -445 -645 125
rect -565 -445 -545 125
rect -465 -445 -445 125
rect -365 -445 -345 125
rect -265 -445 -245 125
rect -165 -445 -145 125
rect -65 -445 -45 125
rect 35 -445 55 125
rect 135 -445 155 125
rect 235 -445 255 125
rect 335 -445 355 125
<< pdiffc >>
rect -665 2640 -645 2760
rect -565 2640 -545 2760
rect -465 2640 -445 2760
rect -365 2640 -345 2760
rect -265 2640 -245 2760
rect -165 2640 -145 2760
rect -65 2640 -45 2760
rect 35 2640 55 2760
rect 135 2640 155 2760
rect 235 2640 255 2760
rect 335 2640 355 2760
rect -665 2140 -645 2410
rect -565 2140 -545 2410
rect -465 2140 -445 2410
rect -365 2140 -345 2410
rect -265 2140 -245 2410
rect -165 2140 -145 2410
rect -65 2140 -45 2410
rect 35 2140 55 2410
rect 135 2140 155 2410
rect 235 2140 255 2410
rect 335 2140 355 2410
rect -665 1265 -645 1835
rect -565 1265 -545 1835
rect -465 1265 -445 1835
rect -365 1265 -345 1835
rect -265 1265 -245 1835
rect -165 1265 -145 1835
rect -65 1265 -45 1835
rect 35 1265 55 1835
rect 135 1265 155 1835
rect 235 1265 255 1835
rect 335 1265 355 1835
<< psubdiff >>
rect -730 125 -680 140
rect -730 -445 -715 125
rect -695 -445 -680 125
rect -730 -460 -680 -445
rect 370 125 420 140
rect 370 -445 385 125
rect 405 -445 420 125
rect 370 -460 420 -445
<< nsubdiff >>
rect -730 2760 -680 2775
rect -730 2640 -715 2760
rect -695 2640 -680 2760
rect -730 2625 -680 2640
rect 370 2760 420 2775
rect 370 2640 385 2760
rect 405 2640 420 2760
rect 370 2625 420 2640
rect -730 2410 -680 2425
rect -730 2140 -715 2410
rect -695 2140 -680 2410
rect -730 2125 -680 2140
rect 370 2410 420 2425
rect 370 2140 385 2410
rect 405 2140 420 2410
rect 370 2125 420 2140
rect -730 1835 -680 1850
rect -730 1265 -715 1835
rect -695 1265 -680 1835
rect -730 1250 -680 1265
rect 370 1835 420 1850
rect 370 1265 385 1835
rect 405 1265 420 1835
rect 370 1250 420 1265
<< psubdiffcont >>
rect -715 -445 -695 125
rect 385 -445 405 125
<< nsubdiffcont >>
rect -715 2640 -695 2760
rect 385 2640 405 2760
rect -715 2140 -695 2410
rect 385 2140 405 2410
rect -715 1265 -695 1835
rect 385 1265 405 1835
<< poly >>
rect -530 2835 -480 2850
rect -530 2810 -520 2835
rect -495 2810 -480 2835
rect -630 2775 -580 2790
rect -530 2775 -480 2810
rect -430 2775 -380 2790
rect -330 2775 -280 2790
rect -230 2775 -180 2790
rect -130 2775 -80 2790
rect -30 2775 20 2790
rect 70 2775 120 2790
rect 170 2775 220 2790
rect 270 2775 320 2790
rect -630 2610 -580 2625
rect -675 2600 -580 2610
rect -675 2580 -665 2600
rect -645 2595 -580 2600
rect -530 2610 -480 2625
rect -430 2610 -380 2625
rect -330 2610 -280 2625
rect -230 2610 -180 2625
rect -130 2610 -80 2625
rect -30 2610 20 2625
rect 70 2610 120 2625
rect 170 2610 220 2625
rect -530 2595 220 2610
rect 270 2610 320 2625
rect 270 2600 365 2610
rect 270 2595 335 2600
rect -645 2580 -635 2595
rect -675 2570 -635 2580
rect 325 2580 335 2595
rect 355 2580 365 2600
rect 325 2570 365 2580
rect 375 2535 415 2545
rect 375 2520 385 2535
rect 105 2515 385 2520
rect 405 2515 415 2535
rect 105 2505 415 2515
rect 105 2480 120 2505
rect -675 2470 -635 2480
rect -675 2450 -665 2470
rect -645 2455 -635 2470
rect -430 2465 120 2480
rect -645 2450 -580 2455
rect -675 2440 -580 2450
rect -630 2425 -580 2440
rect -530 2425 -480 2440
rect -430 2425 -380 2465
rect -330 2425 -280 2465
rect -230 2425 -180 2440
rect -130 2425 -80 2440
rect -30 2425 20 2465
rect 70 2425 120 2465
rect 325 2470 365 2480
rect 325 2455 335 2470
rect 270 2450 335 2455
rect 355 2450 365 2470
rect 270 2440 365 2450
rect 170 2425 220 2440
rect 270 2425 320 2440
rect -630 2110 -580 2125
rect -530 2085 -480 2125
rect -430 2110 -380 2125
rect -330 2110 -280 2125
rect -230 2085 -180 2125
rect -130 2085 -80 2125
rect -30 2110 20 2125
rect 70 2110 120 2125
rect 170 2085 220 2125
rect 270 2110 320 2125
rect -530 2075 325 2085
rect -530 2070 295 2075
rect 285 2055 295 2070
rect 315 2055 325 2075
rect 285 2045 325 2055
rect -375 2035 65 2045
rect -375 2015 -365 2035
rect -345 2030 35 2035
rect -345 2015 -335 2030
rect -375 2005 -335 2015
rect 25 2015 35 2030
rect 55 2015 65 2035
rect 25 2005 65 2015
rect -530 1930 220 1945
rect -675 1895 -635 1905
rect -675 1875 -665 1895
rect -645 1880 -635 1895
rect -645 1875 -580 1880
rect -675 1865 -580 1875
rect -630 1850 -580 1865
rect -530 1850 -480 1930
rect -430 1850 -380 1865
rect -330 1850 -280 1865
rect -230 1850 -180 1930
rect -130 1850 -80 1930
rect -30 1850 20 1865
rect 70 1850 120 1865
rect 170 1850 220 1930
rect 325 1895 365 1905
rect 325 1880 335 1895
rect 270 1875 335 1880
rect 355 1875 365 1895
rect 270 1865 365 1875
rect 270 1850 320 1865
rect -630 1235 -580 1250
rect -725 1210 -685 1220
rect -725 1190 -715 1210
rect -695 1195 -685 1210
rect -530 1195 -480 1250
rect -695 1190 -480 1195
rect -725 1180 -480 1190
rect -430 1210 -380 1250
rect -330 1210 -280 1250
rect -230 1235 -180 1250
rect -130 1235 -80 1250
rect -30 1210 20 1250
rect 70 1210 120 1250
rect 170 1235 220 1250
rect 270 1235 320 1250
rect -430 1200 120 1210
rect -430 1195 -165 1200
rect -430 340 -415 1195
rect -175 1180 -165 1195
rect -145 1195 120 1200
rect -145 1180 -135 1195
rect -175 1170 -135 1180
rect -575 330 -415 340
rect -575 310 -565 330
rect -545 325 -415 330
rect 105 340 120 1195
rect 105 330 265 340
rect 105 325 235 330
rect -545 310 -535 325
rect -575 300 -535 310
rect 225 310 235 325
rect 255 310 265 330
rect 225 300 265 310
rect -725 250 -685 260
rect -725 230 -715 250
rect -695 235 -685 250
rect -695 230 -415 235
rect -725 220 -415 230
rect -430 195 -415 220
rect -675 185 -635 195
rect -675 165 -665 185
rect -645 170 -635 185
rect -430 180 120 195
rect -645 165 -580 170
rect -675 155 -580 165
rect -630 140 -580 155
rect -530 140 -480 155
rect -430 140 -380 180
rect -330 140 -280 180
rect -230 140 -180 155
rect -130 140 -80 155
rect -30 140 20 180
rect 70 140 120 180
rect 325 185 365 195
rect 325 170 335 185
rect 270 165 335 170
rect 355 165 365 185
rect 270 155 365 165
rect 170 140 220 155
rect 270 140 320 155
rect -630 -475 -580 -460
rect -700 -485 -660 -475
rect -700 -505 -690 -485
rect -670 -500 -660 -485
rect -530 -500 -480 -460
rect -430 -475 -380 -460
rect -330 -475 -280 -460
rect -230 -500 -180 -460
rect -130 -500 -80 -460
rect -30 -475 20 -460
rect 70 -475 120 -460
rect 170 -500 220 -460
rect 270 -475 320 -460
rect -670 -505 220 -500
rect -700 -515 220 -505
<< polycont >>
rect -520 2810 -495 2835
rect -665 2580 -645 2600
rect 335 2580 355 2600
rect 385 2515 405 2535
rect -665 2450 -645 2470
rect 335 2450 355 2470
rect 295 2055 315 2075
rect -365 2015 -345 2035
rect 35 2015 55 2035
rect -665 1875 -645 1895
rect 335 1875 355 1895
rect -715 1190 -695 1210
rect -165 1180 -145 1200
rect -565 310 -545 330
rect 235 310 255 330
rect -715 230 -695 250
rect -665 165 -645 185
rect 335 165 355 185
rect -690 -505 -670 -485
<< locali >>
rect -530 2835 -480 2850
rect -530 2820 -520 2835
rect -730 2810 -520 2820
rect -495 2810 -480 2835
rect -730 2800 -480 2810
rect -725 2760 -635 2770
rect -725 2640 -715 2760
rect -695 2640 -665 2760
rect -645 2640 -635 2760
rect -725 2630 -635 2640
rect -575 2760 -535 2770
rect -575 2640 -565 2760
rect -545 2640 -535 2760
rect -575 2630 -535 2640
rect -475 2760 -435 2770
rect -475 2640 -465 2760
rect -445 2640 -435 2760
rect -675 2600 -635 2630
rect -675 2580 -665 2600
rect -645 2580 -635 2600
rect -675 2570 -635 2580
rect -475 2600 -435 2640
rect -375 2760 -335 2770
rect -375 2640 -365 2760
rect -345 2640 -335 2760
rect -375 2630 -335 2640
rect -275 2760 -235 2770
rect -275 2640 -265 2760
rect -245 2640 -235 2760
rect -275 2600 -235 2640
rect -175 2760 -135 2770
rect -175 2640 -165 2760
rect -145 2640 -135 2760
rect -175 2630 -135 2640
rect -75 2760 -35 2770
rect -75 2640 -65 2760
rect -45 2640 -35 2760
rect -75 2600 -35 2640
rect 25 2760 65 2770
rect 25 2640 35 2760
rect 55 2640 65 2760
rect 25 2630 65 2640
rect 125 2760 165 2770
rect 125 2640 135 2760
rect 155 2640 165 2760
rect 125 2600 165 2640
rect 225 2760 265 2770
rect 225 2640 235 2760
rect 255 2640 265 2760
rect 225 2630 265 2640
rect 325 2760 415 2770
rect 325 2640 335 2760
rect 355 2640 385 2760
rect 405 2640 415 2760
rect 325 2630 415 2640
rect -475 2580 165 2600
rect -675 2470 -635 2480
rect -675 2450 -665 2470
rect -645 2450 -635 2470
rect -675 2420 -635 2450
rect -725 2410 -635 2420
rect -725 2140 -715 2410
rect -695 2140 -665 2410
rect -645 2140 -635 2410
rect -725 2130 -635 2140
rect -575 2410 -535 2420
rect -575 2140 -565 2410
rect -545 2140 -535 2410
rect -575 1985 -535 2140
rect -475 2410 -435 2580
rect -475 2140 -465 2410
rect -445 2140 -435 2410
rect -475 2130 -435 2140
rect -375 2410 -335 2420
rect -375 2140 -365 2410
rect -345 2140 -335 2410
rect -375 2045 -335 2140
rect -275 2410 -235 2580
rect -275 2140 -265 2410
rect -245 2140 -235 2410
rect -275 2130 -235 2140
rect -175 2410 -135 2420
rect -175 2140 -165 2410
rect -145 2140 -135 2410
rect -440 2035 -335 2045
rect -440 2015 -430 2035
rect -410 2025 -365 2035
rect -410 2015 -400 2025
rect -440 2005 -400 2015
rect -375 2015 -365 2025
rect -345 2015 -335 2035
rect -375 2005 -335 2015
rect -175 1995 -135 2140
rect -75 2410 -35 2580
rect -75 2140 -65 2410
rect -45 2140 -35 2410
rect -75 2130 -35 2140
rect 25 2410 65 2420
rect 25 2140 35 2410
rect 55 2140 65 2410
rect 25 2035 65 2140
rect 125 2410 165 2580
rect 325 2600 365 2630
rect 325 2580 335 2600
rect 355 2580 365 2600
rect 325 2570 365 2580
rect 375 2535 415 2545
rect 375 2515 385 2535
rect 405 2525 415 2535
rect 405 2515 420 2525
rect 375 2505 420 2515
rect 325 2470 365 2480
rect 325 2450 335 2470
rect 355 2450 365 2470
rect 325 2420 365 2450
rect 125 2140 135 2410
rect 155 2140 165 2410
rect 125 2130 165 2140
rect 225 2410 265 2420
rect 225 2140 235 2410
rect 255 2140 265 2410
rect 25 2015 35 2035
rect 55 2015 65 2035
rect 25 2005 65 2015
rect -175 1985 -165 1995
rect -575 1975 -165 1985
rect -145 1985 -135 1995
rect 225 1985 265 2140
rect 325 2410 415 2420
rect 325 2140 335 2410
rect 355 2140 385 2410
rect 405 2140 415 2410
rect 325 2130 415 2140
rect 285 2075 420 2085
rect 285 2055 295 2075
rect 315 2065 420 2075
rect 315 2055 325 2065
rect 285 2045 325 2055
rect -145 1975 265 1985
rect -575 1965 265 1975
rect -475 1905 165 1925
rect -675 1895 -635 1905
rect -675 1875 -665 1895
rect -645 1875 -635 1895
rect -675 1845 -635 1875
rect -725 1835 -635 1845
rect -725 1265 -715 1835
rect -695 1265 -665 1835
rect -645 1265 -635 1835
rect -725 1255 -635 1265
rect -575 1835 -535 1845
rect -575 1265 -565 1835
rect -545 1265 -535 1835
rect -725 1210 -685 1220
rect -725 1200 -715 1210
rect -730 1190 -715 1200
rect -695 1190 -685 1210
rect -730 1180 -685 1190
rect -575 1150 -535 1265
rect -475 1835 -435 1905
rect -275 1865 -35 1885
rect -475 1265 -465 1835
rect -445 1265 -435 1835
rect -475 1255 -435 1265
rect -375 1835 -335 1845
rect -375 1265 -365 1835
rect -345 1265 -335 1835
rect -375 1255 -335 1265
rect -275 1835 -235 1865
rect -275 1265 -265 1835
rect -245 1265 -235 1835
rect -275 1255 -235 1265
rect -175 1835 -135 1845
rect -175 1265 -165 1835
rect -145 1265 -135 1835
rect -175 1200 -135 1265
rect -75 1835 -35 1865
rect -75 1265 -65 1835
rect -45 1265 -35 1835
rect -75 1255 -35 1265
rect 25 1835 65 1845
rect 25 1265 35 1835
rect 55 1265 65 1835
rect 25 1255 65 1265
rect 125 1835 165 1905
rect 325 1895 365 1905
rect 325 1875 335 1895
rect 355 1875 365 1895
rect 325 1850 365 1875
rect 325 1845 370 1850
rect 125 1265 135 1835
rect 155 1265 165 1835
rect 125 1255 165 1265
rect 225 1835 265 1845
rect 225 1265 235 1835
rect 255 1265 265 1835
rect -175 1180 -165 1200
rect -145 1180 -135 1200
rect -175 1170 -135 1180
rect 225 1150 265 1265
rect 325 1835 415 1845
rect 325 1265 335 1835
rect 355 1265 385 1835
rect 405 1265 415 1835
rect 325 1255 415 1265
rect -575 1130 440 1150
rect -730 1090 -705 1110
rect -725 260 -705 1090
rect -575 330 -535 340
rect -575 310 -565 330
rect -545 310 -535 330
rect -725 250 -685 260
rect -725 230 -715 250
rect -695 230 -685 250
rect -725 220 -685 230
rect -675 185 -635 195
rect -675 165 -665 185
rect -645 165 -635 185
rect -675 140 -635 165
rect -680 135 -635 140
rect -725 125 -635 135
rect -725 -445 -715 125
rect -695 -445 -665 125
rect -645 -445 -635 125
rect -725 -455 -635 -445
rect -575 125 -535 310
rect -575 -445 -565 125
rect -545 -445 -535 125
rect -575 -455 -535 -445
rect -475 290 -435 300
rect -475 270 -465 290
rect -445 270 -435 290
rect -475 125 -435 270
rect -475 -445 -465 125
rect -445 -445 -435 125
rect -700 -485 -660 -475
rect -730 -505 -690 -485
rect -670 -505 -660 -485
rect -700 -515 -660 -505
rect -475 -515 -435 -445
rect -375 125 -335 135
rect -375 -445 -365 125
rect -345 -445 -335 125
rect -375 -455 -335 -445
rect -275 125 -235 135
rect -275 -445 -265 125
rect -245 -445 -235 125
rect -275 -475 -235 -445
rect -175 125 -135 1130
rect 225 330 265 340
rect 225 310 235 330
rect 255 310 265 330
rect -175 -445 -165 125
rect -145 -445 -135 125
rect -175 -455 -135 -445
rect -75 250 -35 260
rect -75 230 -65 250
rect -45 230 -35 250
rect -75 125 -35 230
rect -75 -445 -65 125
rect -45 -445 -35 125
rect -75 -475 -35 -445
rect 25 125 65 135
rect 25 -445 35 125
rect 55 -445 65 125
rect 25 -455 65 -445
rect 125 125 165 135
rect 125 -445 135 125
rect 155 -445 165 125
rect -275 -495 -35 -475
rect 125 -515 165 -445
rect 225 125 265 310
rect 225 -445 235 125
rect 255 -445 265 125
rect 225 -455 265 -445
rect 325 185 365 195
rect 325 165 335 185
rect 355 165 365 185
rect 325 135 365 165
rect 325 125 415 135
rect 325 -445 335 125
rect 355 -445 385 125
rect 405 -445 415 125
rect 325 -455 415 -445
rect -475 -535 165 -515
<< viali >>
rect -715 2640 -695 2760
rect -665 2640 -645 2760
rect -565 2640 -545 2760
rect -365 2640 -345 2760
rect -165 2640 -145 2760
rect 35 2640 55 2760
rect 235 2640 255 2760
rect 335 2640 355 2760
rect 385 2640 405 2760
rect -430 2015 -410 2035
rect -165 1975 -145 1995
rect -715 1265 -695 1835
rect -665 1265 -645 1835
rect -365 1265 -345 1835
rect 35 1265 55 1835
rect 335 1265 355 1835
rect 385 1265 405 1835
rect -715 -445 -695 125
rect -665 -445 -645 125
rect -465 270 -445 290
rect -365 -445 -345 125
rect -65 230 -45 250
rect 35 -445 55 125
rect 335 -445 355 125
rect 385 -445 405 125
<< metal1 >>
rect -730 2760 420 2770
rect -730 2640 -715 2760
rect -695 2640 -665 2760
rect -645 2640 -565 2760
rect -545 2640 -365 2760
rect -345 2640 -165 2760
rect -145 2640 35 2760
rect 55 2640 235 2760
rect 255 2640 335 2760
rect 355 2640 385 2760
rect 405 2640 420 2760
rect -730 2130 420 2640
rect -730 1845 -635 2130
rect -440 2035 -400 2045
rect -440 2015 -430 2035
rect -410 2015 -400 2035
rect -440 1915 -400 2015
rect -175 1995 -135 2005
rect -175 1975 -165 1995
rect -145 1975 -135 1995
rect -175 1915 -135 1975
rect -440 1875 -235 1915
rect -175 1875 -35 1915
rect -730 1835 -335 1845
rect -730 1265 -715 1835
rect -695 1265 -665 1835
rect -645 1265 -365 1835
rect -345 1265 -335 1835
rect -730 1255 -335 1265
rect -275 300 -235 1875
rect -475 290 -235 300
rect -475 270 -465 290
rect -445 270 -235 290
rect -475 260 -235 270
rect -75 250 -35 1875
rect 325 1845 420 2130
rect 25 1835 420 1845
rect 25 1265 35 1835
rect 55 1265 335 1835
rect 355 1265 385 1835
rect 405 1265 420 1835
rect 25 1255 420 1265
rect -75 230 -65 250
rect -45 230 -35 250
rect -75 220 -35 230
rect -725 125 415 135
rect -725 -445 -715 125
rect -695 -445 -665 125
rect -645 -445 -365 125
rect -345 -445 35 125
rect 55 -445 335 125
rect 355 -445 385 125
rect 405 -445 415 125
rect -725 -455 415 -445
<< labels >>
rlabel locali -730 2810 -730 2810 7 Vbp
port 1 w
rlabel metal1 -730 2700 -730 2700 7 VP
port 2 w
rlabel locali -730 1190 -730 1190 7 Vcp
port 3 w
rlabel locali -730 1100 -730 1100 7 Vbn
port 4 w
rlabel psubdiff -730 -165 -730 -165 7 VN
port 5 w
rlabel locali -730 -495 -730 -495 7 Vcn
port 6 w
rlabel locali 440 1140 440 1140 3 Vout
port 7 e
rlabel metal1 420 2075 420 2075 3 V1
port 8 e
rlabel metal1 420 2515 420 2515 3 V2
port 9 e
<< end >>
