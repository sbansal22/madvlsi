magic
tech sky130A
timestamp 1614682669
<< nwell >>
rect -190 655 -20 1240
<< nmos >>
rect -120 300 -105 400
<< pmos >>
rect -120 1000 -105 1095
rect -120 770 -105 865
<< ndiff >>
rect -170 385 -120 400
rect -170 315 -160 385
rect -135 315 -120 385
rect -170 300 -120 315
rect -105 385 -55 400
rect -105 315 -90 385
rect -65 315 -55 385
rect -105 300 -55 315
<< pdiff >>
rect -170 1080 -120 1095
rect -170 1015 -155 1080
rect -135 1015 -120 1080
rect -170 1000 -120 1015
rect -105 1080 -60 1095
rect -105 1015 -90 1080
rect -70 1015 -60 1080
rect -105 1000 -60 1015
rect -170 850 -120 865
rect -170 785 -155 850
rect -135 785 -120 850
rect -170 770 -120 785
rect -105 850 -55 865
rect -105 785 -90 850
rect -70 785 -55 850
rect -105 770 -55 785
<< ndiffc >>
rect -160 315 -135 385
rect -90 315 -65 385
<< pdiffc >>
rect -155 1015 -135 1080
rect -90 1015 -70 1080
rect -155 785 -135 850
rect -90 785 -70 850
<< psubdiff >>
rect -170 125 -120 140
rect -170 55 -155 125
rect -135 55 -120 125
rect -170 40 -120 55
<< nsubdiff >>
rect -170 1205 -120 1220
rect -170 1140 -155 1205
rect -135 1140 -120 1205
rect -170 1125 -120 1140
<< psubdiffcont >>
rect -155 55 -135 125
<< nsubdiffcont >>
rect -155 1140 -135 1205
<< poly >>
rect -120 1095 -105 1110
rect -120 935 -105 1000
rect -165 925 -105 935
rect -165 905 -155 925
rect -135 905 -105 925
rect -165 895 -105 905
rect -120 865 -105 895
rect -120 750 -105 770
rect -165 735 -105 750
rect -165 425 -150 735
rect -120 710 -105 735
rect -120 700 -60 710
rect -120 695 -90 700
rect -100 680 -90 695
rect -70 680 -60 700
rect -100 670 -60 680
rect -165 410 -105 425
rect -120 400 -105 410
rect -120 285 -105 300
<< polycont >>
rect -155 905 -135 925
rect -90 680 -70 700
<< locali >>
rect -165 1205 -125 1215
rect -165 1140 -155 1205
rect -135 1140 -125 1205
rect -165 1130 -125 1140
rect -165 1080 -125 1090
rect -165 1015 -155 1080
rect -135 1015 -125 1080
rect -165 1005 -125 1015
rect -100 1080 -60 1090
rect -100 1015 -90 1080
rect -70 1060 -60 1080
rect -70 1040 -40 1060
rect -70 1015 -60 1040
rect -100 1005 -60 1015
rect -165 925 -125 935
rect -170 905 -155 925
rect -135 905 -125 925
rect -165 895 -125 905
rect -99 860 -80 1005
rect -165 850 -125 860
rect -165 785 -155 850
rect -135 785 -125 850
rect -165 775 -125 785
rect -100 850 -60 860
rect -100 785 -90 850
rect -70 785 -60 850
rect -100 775 -60 785
rect -100 755 -80 775
rect -165 735 -80 755
rect -165 435 -145 735
rect -45 710 -25 735
rect -100 700 -25 710
rect -100 680 -90 700
rect -70 690 -25 700
rect -70 680 -60 690
rect -100 670 -60 680
rect -165 415 -80 435
rect -100 395 -80 415
rect -170 385 -125 395
rect -170 315 -160 385
rect -135 315 -125 385
rect -170 305 -125 315
rect -100 385 -55 395
rect -100 315 -90 385
rect -65 315 -55 385
rect -100 305 -55 315
rect -165 125 -125 135
rect -165 55 -155 125
rect -135 55 -125 125
rect -165 45 -125 55
rect -190 5 -45 25
<< viali >>
rect -155 1140 -135 1205
rect -155 1015 -135 1080
rect -155 785 -135 850
rect -160 315 -135 385
rect -155 55 -135 125
<< metal1 >>
rect -170 1205 -45 1220
rect -170 1140 -155 1205
rect -135 1140 -45 1205
rect -170 1125 -45 1140
rect -170 1080 -125 1125
rect -170 1015 -155 1080
rect -135 1015 -125 1080
rect -170 850 -125 1015
rect -170 785 -155 850
rect -135 785 -125 850
rect -170 770 -125 785
rect -170 385 -125 400
rect -170 315 -160 385
rect -135 315 -125 385
rect -170 140 -125 315
rect -170 125 -45 140
rect -170 55 -155 125
rect -135 55 -45 125
rect -170 40 -45 55
<< labels >>
rlabel metal1 -170 1170 -170 1170 7 VP
port 1 w
rlabel locali -170 915 -170 915 7 D
port 2 w
rlabel metal1 -170 90 -170 90 7 VN
port 3 w
rlabel locali -190 15 -190 15 7 CLK
port 4 w
rlabel locali -25 720 -25 720 3 D
port 5 e
rlabel locali -40 1050 -40 1050 3 Dn
port 6 e
<< end >>
