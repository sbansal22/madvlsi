magic
tech sky130A
timestamp 1614269894
<< nmos >>
rect 0 420 15 620
rect 65 520 80 620
rect 130 520 145 620
rect 195 520 210 620
rect 0 -5 15 195
rect 65 -5 80 95
rect 130 -5 145 95
rect 195 -5 210 95
<< ndiff >>
rect -50 605 0 620
rect -50 535 -35 605
rect -15 535 0 605
rect -50 420 0 535
rect 15 520 65 620
rect 80 605 130 620
rect 80 535 95 605
rect 115 535 130 605
rect 80 520 130 535
rect 145 605 195 620
rect 145 535 160 605
rect 180 535 195 605
rect 145 520 195 535
rect 210 605 260 620
rect 210 535 225 605
rect 245 535 260 605
rect 210 520 260 535
rect 15 420 50 520
rect -50 80 0 195
rect -50 10 -35 80
rect -15 10 0 80
rect -50 -5 0 10
rect 15 95 50 195
rect 15 -5 65 95
rect 80 80 130 95
rect 80 10 95 80
rect 115 10 130 80
rect 80 -5 130 10
rect 145 80 195 95
rect 145 10 160 80
rect 180 10 195 80
rect 145 -5 195 10
rect 210 80 255 95
rect 210 10 225 80
rect 245 10 255 80
rect 210 -5 255 10
<< ndiffc >>
rect -35 535 -15 605
rect 95 535 115 605
rect 160 535 180 605
rect 225 535 245 605
rect -35 10 -15 80
rect 95 10 115 80
rect 160 10 180 80
rect 225 10 245 80
<< psubdiff >>
rect -100 605 -50 620
rect -100 535 -85 605
rect -65 535 -50 605
rect -100 420 -50 535
rect 260 605 310 620
rect 260 535 275 605
rect 295 535 310 605
rect 260 520 310 535
rect -100 80 -50 195
rect -100 10 -85 80
rect -60 10 -50 80
rect -100 -5 -50 10
rect 255 80 305 95
rect 255 10 265 80
rect 290 10 305 80
rect 255 -5 305 10
<< psubdiffcont >>
rect -85 535 -65 605
rect 275 535 295 605
rect -85 10 -60 80
rect 265 10 290 80
<< poly >>
rect 0 620 15 710
rect 65 620 80 710
rect 130 620 145 710
rect 195 620 210 710
rect 0 195 15 420
rect 65 410 80 520
rect 40 400 80 410
rect 40 380 50 400
rect 70 380 80 400
rect 40 370 80 380
rect 65 335 105 345
rect 65 315 75 335
rect 95 315 105 335
rect 65 305 105 315
rect 65 95 80 305
rect 130 95 145 520
rect 195 510 210 520
rect 170 495 210 510
rect 170 185 185 495
rect 210 460 250 470
rect 210 440 220 460
rect 240 440 250 460
rect 210 430 250 440
rect 170 175 210 185
rect 170 155 180 175
rect 200 155 210 175
rect 170 145 210 155
rect 235 120 250 430
rect 195 105 250 120
rect 195 95 210 105
rect 0 -20 15 -5
rect -25 -30 15 -20
rect -25 -50 -15 -30
rect 5 -50 15 -30
rect -25 -60 15 -50
rect 65 -55 80 -5
rect 130 -20 145 -5
rect 105 -30 145 -20
rect 105 -50 115 -30
rect 135 -50 145 -30
rect 105 -60 145 -50
rect 195 -55 210 -5
<< polycont >>
rect 50 380 70 400
rect 75 315 95 335
rect 220 440 240 460
rect 180 155 200 175
rect -15 -50 5 -30
rect 115 -50 135 -30
<< locali >>
rect -95 605 -5 615
rect -95 535 -85 605
rect -65 535 -35 605
rect -15 535 -5 605
rect -95 525 -5 535
rect 85 605 125 615
rect 85 535 95 605
rect 115 535 125 605
rect 85 525 125 535
rect 150 605 190 615
rect 150 535 160 605
rect 180 535 190 605
rect 150 525 190 535
rect 215 605 305 615
rect 215 535 225 605
rect 245 535 275 605
rect 295 535 305 605
rect 215 525 305 535
rect 40 400 80 410
rect 40 390 50 400
rect 20 380 50 390
rect 70 380 80 400
rect 20 370 80 380
rect 20 90 40 370
rect 105 345 125 525
rect 170 470 190 525
rect 170 460 250 470
rect 170 450 220 460
rect 210 440 220 450
rect 240 440 250 460
rect 210 430 250 440
rect 65 335 125 345
rect 65 315 75 335
rect 95 325 125 335
rect 95 315 105 325
rect 65 305 105 315
rect 170 175 210 185
rect 170 155 180 175
rect 200 155 210 175
rect 170 145 210 155
rect 170 90 190 145
rect -95 80 -5 90
rect -95 10 -85 80
rect -60 10 -35 80
rect -15 10 -5 80
rect 20 80 125 90
rect 20 70 95 80
rect -95 0 -5 10
rect 85 10 95 70
rect 115 10 125 80
rect 85 0 125 10
rect 150 80 190 90
rect 150 10 160 80
rect 180 10 190 80
rect 150 0 190 10
rect 215 80 300 90
rect 215 10 225 80
rect 245 10 265 80
rect 290 10 300 80
rect 215 0 300 10
rect -120 -30 280 -20
rect -120 -40 -15 -30
rect -25 -50 -15 -40
rect 5 -40 115 -30
rect 5 -50 15 -40
rect -25 -60 15 -50
rect 105 -50 115 -40
rect 135 -40 280 -30
rect 135 -50 145 -40
rect 105 -60 145 -50
<< viali >>
rect -85 535 -65 605
rect 275 535 295 605
rect -85 10 -60 80
rect 265 10 290 80
<< metal1 >>
rect -115 605 330 615
rect -115 535 -85 605
rect -65 535 275 605
rect 295 535 330 605
rect -115 525 330 535
rect -120 80 325 90
rect -120 10 -85 80
rect -60 10 265 80
rect 290 10 325 80
rect -120 0 325 10
<< end >>
