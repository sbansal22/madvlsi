magic
tech sky130A
timestamp 1613291521
<< nwell >>
rect -120 65 150 220
<< nmos >>
rect 0 -70 15 30
rect 65 -70 80 30
<< pmos >>
rect 0 95 15 195
rect 65 95 80 195
<< ndiff >>
rect -50 15 0 30
rect -50 -55 -35 15
rect -15 -55 0 15
rect -50 -70 0 -55
rect 15 -70 65 30
rect 80 15 130 30
rect 80 -55 95 15
rect 115 -55 130 15
rect 80 -70 130 -55
<< pdiff >>
rect -50 180 0 195
rect -50 110 -35 180
rect -15 110 0 180
rect -50 95 0 110
rect 15 180 65 195
rect 15 110 30 180
rect 50 110 65 180
rect 15 95 65 110
rect 80 180 130 195
rect 80 110 95 180
rect 115 110 130 180
rect 80 95 130 110
<< ndiffc >>
rect -35 -55 -15 15
rect 95 -55 115 15
<< pdiffc >>
rect -35 110 -15 180
rect 30 110 50 180
rect 95 110 115 180
<< psubdiff >>
rect -100 15 -50 30
rect -100 -55 -85 15
rect -65 -55 -50 15
rect -100 -70 -50 -55
<< nsubdiff >>
rect -100 180 -50 195
rect -100 110 -85 180
rect -65 110 -50 180
rect -100 95 -50 110
<< psubdiffcont >>
rect -85 -55 -65 15
<< nsubdiffcont >>
rect -85 110 -65 180
<< poly >>
rect 0 195 15 220
rect 65 195 80 220
rect 0 30 15 95
rect 65 30 80 95
rect 0 -85 15 -70
rect -25 -95 15 -85
rect -25 -115 -15 -95
rect 5 -115 15 -95
rect -25 -125 15 -115
rect 65 -150 80 -70
rect 40 -160 80 -150
rect 40 -180 50 -160
rect 70 -180 80 -160
rect 40 -190 80 -180
<< polycont >>
rect -15 -115 5 -95
rect 50 -180 70 -160
<< locali >>
rect -95 180 -5 190
rect -95 110 -85 180
rect -65 110 -35 180
rect -15 110 -5 180
rect -95 100 -5 110
rect 20 180 60 190
rect 20 110 30 180
rect 50 110 60 180
rect 20 100 60 110
rect 85 180 125 190
rect 85 110 95 180
rect 115 110 125 180
rect 85 100 125 110
rect 40 25 60 100
rect -95 15 -5 25
rect -95 -55 -85 15
rect -65 -55 -35 15
rect -15 -55 -5 15
rect 40 15 125 25
rect 40 5 95 15
rect -95 -65 -5 -55
rect 85 -55 95 5
rect 115 -55 125 15
rect 85 -65 125 -55
rect 105 -85 125 -65
rect -120 -95 15 -85
rect -120 -105 -15 -95
rect -25 -115 -15 -105
rect 5 -115 15 -95
rect 105 -105 150 -85
rect -25 -125 15 -115
rect -120 -160 80 -150
rect -120 -170 50 -160
rect 40 -180 50 -170
rect 70 -180 80 -160
rect 40 -190 80 -180
<< viali >>
rect -85 110 -65 180
rect -35 110 -15 180
rect 95 110 115 180
rect -85 -55 -65 15
rect -35 -55 -15 15
<< metal1 >>
rect -120 180 150 190
rect -120 110 -85 180
rect -65 110 -35 180
rect -15 110 95 180
rect 115 110 150 180
rect -120 100 150 110
rect -120 15 150 25
rect -120 -55 -85 15
rect -65 -55 -35 15
rect -15 -55 150 15
rect -120 -65 150 -55
<< labels >>
rlabel metal1 -120 145 -120 145 7 VP
port 4 w
rlabel locali 150 -95 150 -95 3 Y
port 2 e
rlabel locali -120 -160 -120 -160 7 B
port 3 w
rlabel locali -120 -95 -120 -95 7 A
port 1 w
rlabel metal1 -120 -20 -120 -20 7 VN
port 5 w
<< end >>
