magic
tech sky130A
timestamp 1615670771
<< nwell >>
rect -70 3680 1320 4320
rect -70 2430 1320 3070
<< nmos >>
rect 50 1200 100 1800
rect 150 1200 200 1800
rect 250 1200 300 1800
rect 350 1200 400 1800
rect 550 1200 600 1800
rect 650 1200 700 1800
rect 850 1200 900 1800
rect 950 1200 1000 1800
rect 1050 1200 1100 1800
rect 1150 1200 1200 1800
rect 50 0 100 600
rect 150 0 200 600
rect 250 0 300 600
rect 350 0 400 600
rect 550 0 600 600
rect 650 0 700 600
rect 850 0 900 600
rect 950 0 1000 600
rect 1050 0 1100 600
rect 1150 0 1200 600
<< pmos >>
rect 50 3700 100 4300
rect 150 3700 200 4300
rect 250 3700 300 4300
rect 350 3700 400 4300
rect 550 3700 600 4300
rect 650 3700 700 4300
rect 850 3700 900 4300
rect 950 3700 1000 4300
rect 1050 3700 1100 4300
rect 1150 3700 1200 4300
rect 50 2450 100 3050
rect 150 2450 200 3050
rect 250 2450 300 3050
rect 350 2450 400 3050
rect 550 2450 600 3050
rect 650 2450 700 3050
rect 850 2450 900 3050
rect 950 2450 1000 3050
rect 1050 2450 1100 3050
rect 1150 2450 1200 3050
<< ndiff >>
rect 0 1785 50 1800
rect 0 1215 15 1785
rect 35 1215 50 1785
rect 0 1200 50 1215
rect 100 1785 150 1800
rect 100 1215 115 1785
rect 135 1215 150 1785
rect 100 1200 150 1215
rect 200 1785 250 1800
rect 200 1215 215 1785
rect 235 1215 250 1785
rect 200 1200 250 1215
rect 300 1785 350 1800
rect 300 1215 315 1785
rect 335 1215 350 1785
rect 300 1200 350 1215
rect 400 1785 450 1800
rect 400 1215 415 1785
rect 435 1215 450 1785
rect 400 1200 450 1215
rect 500 1785 550 1800
rect 500 1215 515 1785
rect 535 1215 550 1785
rect 500 1200 550 1215
rect 600 1785 650 1800
rect 600 1215 615 1785
rect 635 1215 650 1785
rect 600 1200 650 1215
rect 700 1785 750 1800
rect 700 1215 715 1785
rect 735 1215 750 1785
rect 700 1200 750 1215
rect 800 1785 850 1800
rect 800 1215 815 1785
rect 835 1215 850 1785
rect 800 1200 850 1215
rect 900 1785 950 1800
rect 900 1215 915 1785
rect 935 1215 950 1785
rect 900 1200 950 1215
rect 1000 1785 1050 1800
rect 1000 1215 1015 1785
rect 1035 1215 1050 1785
rect 1000 1200 1050 1215
rect 1100 1785 1150 1800
rect 1100 1215 1115 1785
rect 1135 1215 1150 1785
rect 1100 1200 1150 1215
rect 1200 1785 1250 1800
rect 1200 1215 1215 1785
rect 1235 1215 1250 1785
rect 1200 1200 1250 1215
rect 0 585 50 600
rect 0 15 15 585
rect 35 15 50 585
rect 0 0 50 15
rect 100 585 150 600
rect 100 15 115 585
rect 135 15 150 585
rect 100 0 150 15
rect 200 585 250 600
rect 200 15 215 585
rect 235 15 250 585
rect 200 0 250 15
rect 300 585 350 600
rect 300 15 315 585
rect 335 15 350 585
rect 300 0 350 15
rect 400 585 450 600
rect 400 15 415 585
rect 435 15 450 585
rect 400 0 450 15
rect 500 585 550 600
rect 500 15 515 585
rect 535 15 550 585
rect 500 0 550 15
rect 600 585 650 600
rect 600 15 615 585
rect 635 15 650 585
rect 600 0 650 15
rect 700 585 750 600
rect 700 15 715 585
rect 735 15 750 585
rect 700 0 750 15
rect 800 585 850 600
rect 800 15 815 585
rect 835 15 850 585
rect 800 0 850 15
rect 900 585 950 600
rect 900 15 915 585
rect 935 15 950 585
rect 900 0 950 15
rect 1000 585 1050 600
rect 1000 15 1015 585
rect 1035 15 1050 585
rect 1000 0 1050 15
rect 1100 585 1150 600
rect 1100 15 1115 585
rect 1135 15 1150 585
rect 1100 0 1150 15
rect 1200 585 1250 600
rect 1200 15 1215 585
rect 1235 15 1250 585
rect 1200 0 1250 15
<< pdiff >>
rect 0 4285 50 4300
rect 0 3715 15 4285
rect 35 3715 50 4285
rect 0 3700 50 3715
rect 100 4285 150 4300
rect 100 3715 115 4285
rect 135 3715 150 4285
rect 100 3700 150 3715
rect 200 4285 250 4300
rect 200 3715 215 4285
rect 235 3715 250 4285
rect 200 3700 250 3715
rect 300 4285 350 4300
rect 300 3715 315 4285
rect 335 3715 350 4285
rect 300 3700 350 3715
rect 400 4285 450 4300
rect 400 3715 415 4285
rect 435 3715 450 4285
rect 400 3700 450 3715
rect 500 4285 550 4300
rect 500 3715 515 4285
rect 535 3715 550 4285
rect 500 3700 550 3715
rect 600 4285 650 4300
rect 600 3715 615 4285
rect 635 3715 650 4285
rect 600 3700 650 3715
rect 700 4285 750 4300
rect 700 3715 715 4285
rect 735 3715 750 4285
rect 700 3700 750 3715
rect 800 4285 850 4300
rect 800 3715 815 4285
rect 835 3715 850 4285
rect 800 3700 850 3715
rect 900 4285 950 4300
rect 900 3715 915 4285
rect 935 3715 950 4285
rect 900 3700 950 3715
rect 1000 4285 1050 4300
rect 1000 3715 1015 4285
rect 1035 3715 1050 4285
rect 1000 3700 1050 3715
rect 1100 4285 1150 4300
rect 1100 3715 1115 4285
rect 1135 3715 1150 4285
rect 1100 3700 1150 3715
rect 1200 4285 1250 4300
rect 1200 3715 1215 4285
rect 1235 3715 1250 4285
rect 1200 3700 1250 3715
rect 0 3035 50 3050
rect 0 2465 15 3035
rect 35 2465 50 3035
rect 0 2450 50 2465
rect 100 3035 150 3050
rect 100 2465 115 3035
rect 135 2465 150 3035
rect 100 2450 150 2465
rect 200 3035 250 3050
rect 200 2465 215 3035
rect 235 2465 250 3035
rect 200 2450 250 2465
rect 300 3035 350 3050
rect 300 2465 315 3035
rect 335 2465 350 3035
rect 300 2450 350 2465
rect 400 3035 450 3050
rect 400 2465 415 3035
rect 435 2465 450 3035
rect 400 2450 450 2465
rect 500 3035 550 3050
rect 500 2465 515 3035
rect 535 2465 550 3035
rect 500 2450 550 2465
rect 600 3035 650 3050
rect 600 2465 615 3035
rect 635 2465 650 3035
rect 600 2450 650 2465
rect 700 3035 750 3050
rect 700 2465 715 3035
rect 735 2465 750 3035
rect 700 2450 750 2465
rect 800 3035 850 3050
rect 800 2465 815 3035
rect 835 2465 850 3035
rect 800 2450 850 2465
rect 900 3035 950 3050
rect 900 2465 915 3035
rect 935 2465 950 3035
rect 900 2450 950 2465
rect 1000 3035 1050 3050
rect 1000 2465 1015 3035
rect 1035 2465 1050 3035
rect 1000 2450 1050 2465
rect 1100 3035 1150 3050
rect 1100 2465 1115 3035
rect 1135 2465 1150 3035
rect 1100 2450 1150 2465
rect 1200 3035 1250 3050
rect 1200 2465 1215 3035
rect 1235 2465 1250 3035
rect 1200 2450 1250 2465
<< ndiffc >>
rect 15 1215 35 1785
rect 115 1215 135 1785
rect 215 1215 235 1785
rect 315 1215 335 1785
rect 415 1215 435 1785
rect 515 1215 535 1785
rect 615 1215 635 1785
rect 715 1215 735 1785
rect 815 1215 835 1785
rect 915 1215 935 1785
rect 1015 1215 1035 1785
rect 1115 1215 1135 1785
rect 1215 1215 1235 1785
rect 15 15 35 585
rect 115 15 135 585
rect 215 15 235 585
rect 315 15 335 585
rect 415 15 435 585
rect 515 15 535 585
rect 615 15 635 585
rect 715 15 735 585
rect 815 15 835 585
rect 915 15 935 585
rect 1015 15 1035 585
rect 1115 15 1135 585
rect 1215 15 1235 585
<< pdiffc >>
rect 15 3715 35 4285
rect 115 3715 135 4285
rect 215 3715 235 4285
rect 315 3715 335 4285
rect 415 3715 435 4285
rect 515 3715 535 4285
rect 615 3715 635 4285
rect 715 3715 735 4285
rect 815 3715 835 4285
rect 915 3715 935 4285
rect 1015 3715 1035 4285
rect 1115 3715 1135 4285
rect 1215 3715 1235 4285
rect 15 2465 35 3035
rect 115 2465 135 3035
rect 215 2465 235 3035
rect 315 2465 335 3035
rect 415 2465 435 3035
rect 515 2465 535 3035
rect 615 2465 635 3035
rect 715 2465 735 3035
rect 815 2465 835 3035
rect 915 2465 935 3035
rect 1015 2465 1035 3035
rect 1115 2465 1135 3035
rect 1215 2465 1235 3035
<< psubdiff >>
rect -50 1785 0 1800
rect -50 1215 -35 1785
rect -15 1215 0 1785
rect -50 1200 0 1215
rect 1250 1785 1300 1800
rect 1250 1215 1265 1785
rect 1285 1215 1300 1785
rect 1250 1200 1300 1215
rect -50 585 0 600
rect -50 15 -35 585
rect -15 15 0 585
rect -50 0 0 15
rect 1250 585 1300 600
rect 1250 15 1265 585
rect 1285 15 1300 585
rect 1250 0 1300 15
<< nsubdiff >>
rect -50 4285 0 4300
rect -50 3715 -35 4285
rect -15 3715 0 4285
rect -50 3700 0 3715
rect 1250 4285 1300 4300
rect 1250 3715 1265 4285
rect 1285 3715 1300 4285
rect 1250 3700 1300 3715
rect -50 3035 0 3050
rect -50 2465 -35 3035
rect -15 2465 0 3035
rect -50 2450 0 2465
rect 1250 3035 1300 3050
rect 1250 2465 1265 3035
rect 1285 2465 1300 3035
rect 1250 2450 1300 2465
<< psubdiffcont >>
rect -35 1215 -15 1785
rect 1265 1215 1285 1785
rect -35 15 -15 585
rect 1265 15 1285 585
<< nsubdiffcont >>
rect -35 3715 -15 4285
rect 1265 3715 1285 4285
rect -35 2465 -15 3035
rect 1265 2465 1285 3035
<< poly >>
rect 50 4300 100 4315
rect 150 4300 200 4315
rect 250 4300 300 4315
rect 350 4300 400 4315
rect 550 4300 600 4315
rect 650 4300 700 4315
rect 850 4300 900 4315
rect 950 4300 1000 4315
rect 1050 4300 1100 4315
rect 1150 4300 1200 4315
rect 50 3685 100 3700
rect 150 3685 200 3700
rect 250 3685 300 3700
rect 350 3685 400 3700
rect 550 3685 600 3700
rect 650 3685 700 3700
rect 850 3685 900 3700
rect 950 3685 1000 3700
rect 1050 3685 1100 3700
rect 1150 3685 1200 3700
rect 50 3050 100 3065
rect 150 3050 200 3065
rect 250 3050 300 3065
rect 350 3050 400 3065
rect 550 3050 600 3065
rect 650 3050 700 3065
rect 850 3050 900 3065
rect 950 3050 1000 3065
rect 1050 3050 1100 3065
rect 1150 3050 1200 3065
rect 50 2435 100 2450
rect 150 2435 200 2450
rect 250 2435 300 2450
rect 350 2435 400 2450
rect 550 2435 600 2450
rect 650 2435 700 2450
rect 850 2435 900 2450
rect 950 2435 1000 2450
rect 1050 2435 1100 2450
rect 1150 2435 1200 2450
rect 50 1800 100 1815
rect 150 1800 200 1815
rect 250 1800 300 1815
rect 350 1800 400 1815
rect 550 1800 600 1815
rect 650 1800 700 1815
rect 850 1800 900 1815
rect 950 1800 1000 1815
rect 1050 1800 1100 1815
rect 1150 1800 1200 1815
rect 50 1185 100 1200
rect 150 1185 200 1200
rect 250 1185 300 1200
rect 350 1185 400 1200
rect 550 1185 600 1200
rect 650 1185 700 1200
rect 850 1185 900 1200
rect 950 1185 1000 1200
rect 1050 1185 1100 1200
rect 1150 1185 1200 1200
rect 50 600 100 615
rect 150 600 200 615
rect 250 600 300 615
rect 350 600 400 615
rect 550 600 600 615
rect 650 600 700 615
rect 850 600 900 615
rect 950 600 1000 615
rect 1050 600 1100 615
rect 1150 600 1200 615
rect 50 -15 100 0
rect 150 -15 200 0
rect 250 -15 300 0
rect 350 -15 400 0
rect 550 -15 600 0
rect 650 -15 700 0
rect 850 -15 900 0
rect 950 -15 1000 0
rect 1050 -15 1100 0
rect 1150 -15 1200 0
<< locali >>
rect -45 4285 45 4295
rect -45 3715 -35 4285
rect -15 3715 15 4285
rect 35 3715 45 4285
rect -45 3705 45 3715
rect 105 4285 145 4295
rect 105 3715 115 4285
rect 135 3715 145 4285
rect 105 3705 145 3715
rect 205 4285 245 4295
rect 205 3715 215 4285
rect 235 3715 245 4285
rect 205 3705 245 3715
rect 305 4285 345 4295
rect 305 3715 315 4285
rect 335 3715 345 4285
rect 305 3705 345 3715
rect 405 4285 445 4295
rect 405 3715 415 4285
rect 435 3715 445 4285
rect 405 3705 445 3715
rect 505 4285 545 4295
rect 505 3715 515 4285
rect 535 3715 545 4285
rect 505 3705 545 3715
rect 605 4285 645 4295
rect 605 3715 615 4285
rect 635 3715 645 4285
rect 605 3705 645 3715
rect 705 4285 745 4295
rect 705 3715 715 4285
rect 735 3715 745 4285
rect 705 3705 745 3715
rect 805 4285 845 4295
rect 805 3715 815 4285
rect 835 3715 845 4285
rect 805 3705 845 3715
rect 905 4285 945 4295
rect 905 3715 915 4285
rect 935 3715 945 4285
rect 905 3705 945 3715
rect 1005 4285 1045 4295
rect 1005 3715 1015 4285
rect 1035 3715 1045 4285
rect 1005 3705 1045 3715
rect 1105 4285 1145 4295
rect 1105 3715 1115 4285
rect 1135 3715 1145 4285
rect 1105 3705 1145 3715
rect 1205 4285 1295 4295
rect 1205 3715 1215 4285
rect 1235 3715 1265 4285
rect 1285 3715 1295 4285
rect 1205 3705 1295 3715
rect -45 3035 45 3045
rect -45 2465 -35 3035
rect -15 2465 15 3035
rect 35 2465 45 3035
rect -45 2455 45 2465
rect 105 3035 145 3045
rect 105 2465 115 3035
rect 135 2465 145 3035
rect 105 2455 145 2465
rect 205 3035 245 3045
rect 205 2465 215 3035
rect 235 2465 245 3035
rect 205 2455 245 2465
rect 305 3035 345 3045
rect 305 2465 315 3035
rect 335 2465 345 3035
rect 305 2455 345 2465
rect 405 3035 445 3045
rect 405 2465 415 3035
rect 435 2465 445 3035
rect 405 2455 445 2465
rect 505 3035 545 3045
rect 505 2465 515 3035
rect 535 2465 545 3035
rect 505 2455 545 2465
rect 605 3035 645 3045
rect 605 2465 615 3035
rect 635 2465 645 3035
rect 605 2455 645 2465
rect 705 3035 745 3045
rect 705 2465 715 3035
rect 735 2465 745 3035
rect 705 2455 745 2465
rect 805 3035 845 3045
rect 805 2465 815 3035
rect 835 2465 845 3035
rect 805 2455 845 2465
rect 905 3035 945 3045
rect 905 2465 915 3035
rect 935 2465 945 3035
rect 905 2455 945 2465
rect 1005 3035 1045 3045
rect 1005 2465 1015 3035
rect 1035 2465 1045 3035
rect 1005 2455 1045 2465
rect 1105 3035 1145 3045
rect 1105 2465 1115 3035
rect 1135 2465 1145 3035
rect 1105 2455 1145 2465
rect 1205 3035 1295 3045
rect 1205 2465 1215 3035
rect 1235 2465 1265 3035
rect 1285 2465 1295 3035
rect 1205 2455 1295 2465
rect -45 1785 45 1795
rect -45 1215 -35 1785
rect -15 1215 15 1785
rect 35 1215 45 1785
rect -45 1205 45 1215
rect 105 1785 145 1795
rect 105 1215 115 1785
rect 135 1215 145 1785
rect 105 1205 145 1215
rect 205 1785 245 1795
rect 205 1215 215 1785
rect 235 1215 245 1785
rect 205 1205 245 1215
rect 305 1785 345 1795
rect 305 1215 315 1785
rect 335 1215 345 1785
rect 305 1205 345 1215
rect 405 1785 445 1795
rect 405 1215 415 1785
rect 435 1215 445 1785
rect 405 1205 445 1215
rect 505 1785 545 1795
rect 505 1215 515 1785
rect 535 1215 545 1785
rect 505 1205 545 1215
rect 605 1785 645 1795
rect 605 1215 615 1785
rect 635 1215 645 1785
rect 605 1205 645 1215
rect 705 1785 745 1795
rect 705 1215 715 1785
rect 735 1215 745 1785
rect 705 1205 745 1215
rect 805 1785 845 1795
rect 805 1215 815 1785
rect 835 1215 845 1785
rect 805 1205 845 1215
rect 905 1785 945 1795
rect 905 1215 915 1785
rect 935 1215 945 1785
rect 905 1205 945 1215
rect 1005 1785 1045 1795
rect 1005 1215 1015 1785
rect 1035 1215 1045 1785
rect 1005 1205 1045 1215
rect 1105 1785 1145 1795
rect 1105 1215 1115 1785
rect 1135 1215 1145 1785
rect 1105 1205 1145 1215
rect 1205 1785 1295 1795
rect 1205 1215 1215 1785
rect 1235 1215 1265 1785
rect 1285 1215 1295 1785
rect 1205 1205 1295 1215
rect -45 585 45 595
rect -45 15 -35 585
rect -15 15 15 585
rect 35 15 45 585
rect -45 5 45 15
rect 105 585 145 595
rect 105 15 115 585
rect 135 15 145 585
rect 105 5 145 15
rect 205 585 245 595
rect 205 15 215 585
rect 235 15 245 585
rect 205 5 245 15
rect 305 585 345 595
rect 305 15 315 585
rect 335 15 345 585
rect 305 5 345 15
rect 405 585 445 595
rect 405 15 415 585
rect 435 15 445 585
rect 405 5 445 15
rect 505 585 545 595
rect 505 15 515 585
rect 535 15 545 585
rect 505 5 545 15
rect 605 585 645 595
rect 605 15 615 585
rect 635 15 645 585
rect 605 5 645 15
rect 705 585 745 595
rect 705 15 715 585
rect 735 15 745 585
rect 705 5 745 15
rect 805 585 845 595
rect 805 15 815 585
rect 835 15 845 585
rect 805 5 845 15
rect 905 585 945 595
rect 905 15 915 585
rect 935 15 945 585
rect 905 5 945 15
rect 1005 585 1045 595
rect 1005 15 1015 585
rect 1035 15 1045 585
rect 1005 5 1045 15
rect 1105 585 1145 595
rect 1105 15 1115 585
rect 1135 15 1145 585
rect 1105 5 1145 15
rect 1205 585 1295 595
rect 1205 15 1215 585
rect 1235 15 1265 585
rect 1285 15 1295 585
rect 1205 5 1295 15
<< end >>
