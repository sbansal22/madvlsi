magic
tech sky130A
timestamp 1615805148
<< nwell >>
rect -750 1245 440 3620
<< nmos >>
rect -630 15 -580 615
rect -530 15 -480 615
rect -430 15 -380 615
rect -330 15 -280 615
rect -230 15 -180 615
rect -130 15 -80 615
rect -30 15 20 615
rect 70 15 120 615
rect 170 15 220 615
rect 270 15 320 615
<< pmos >>
rect -630 3465 -580 3600
rect -530 3465 -480 3600
rect -430 3465 -380 3600
rect -330 3465 -280 3600
rect -230 3465 -180 3600
rect -130 3465 -80 3600
rect -30 3465 20 3600
rect 70 3465 120 3600
rect 170 3465 220 3600
rect 270 3465 320 3600
rect -630 2515 -580 2815
rect -530 2515 -480 2815
rect -430 2515 -380 2815
rect -330 2515 -280 2815
rect -230 2515 -180 2815
rect -130 2515 -80 2815
rect -30 2515 20 2815
rect 70 2515 120 2815
rect 170 2515 220 2815
rect 270 2515 320 2815
rect -630 1265 -580 1865
rect -530 1265 -480 1865
rect -430 1265 -380 1865
rect -330 1265 -280 1865
rect -230 1265 -180 1865
rect -130 1265 -80 1865
rect -30 1265 20 1865
rect 70 1265 120 1865
rect 170 1265 220 1865
rect 270 1265 320 1865
<< ndiff >>
rect -680 600 -630 615
rect -680 30 -665 600
rect -645 30 -630 600
rect -680 15 -630 30
rect -580 600 -530 615
rect -580 30 -565 600
rect -545 30 -530 600
rect -580 15 -530 30
rect -480 600 -430 615
rect -480 30 -465 600
rect -445 30 -430 600
rect -480 15 -430 30
rect -380 600 -330 615
rect -380 30 -365 600
rect -345 30 -330 600
rect -380 15 -330 30
rect -280 600 -230 615
rect -280 30 -265 600
rect -245 30 -230 600
rect -280 15 -230 30
rect -180 600 -130 615
rect -180 30 -165 600
rect -145 30 -130 600
rect -180 15 -130 30
rect -80 600 -30 615
rect -80 30 -65 600
rect -45 30 -30 600
rect -80 15 -30 30
rect 20 600 70 615
rect 20 30 35 600
rect 55 30 70 600
rect 20 15 70 30
rect 120 600 170 615
rect 120 30 135 600
rect 155 30 170 600
rect 120 15 170 30
rect 220 600 270 615
rect 220 30 235 600
rect 255 30 270 600
rect 220 15 270 30
rect 320 600 370 615
rect 320 30 335 600
rect 355 30 370 600
rect 320 15 370 30
<< pdiff >>
rect -680 3585 -630 3600
rect -680 3480 -665 3585
rect -645 3480 -630 3585
rect -680 3465 -630 3480
rect -580 3585 -530 3600
rect -580 3480 -565 3585
rect -545 3480 -530 3585
rect -580 3465 -530 3480
rect -480 3585 -430 3600
rect -480 3480 -465 3585
rect -445 3480 -430 3585
rect -480 3465 -430 3480
rect -380 3585 -330 3600
rect -380 3480 -365 3585
rect -345 3480 -330 3585
rect -380 3465 -330 3480
rect -280 3585 -230 3600
rect -280 3480 -265 3585
rect -245 3480 -230 3585
rect -280 3465 -230 3480
rect -180 3585 -130 3600
rect -180 3480 -165 3585
rect -145 3480 -130 3585
rect -180 3465 -130 3480
rect -80 3585 -30 3600
rect -80 3480 -65 3585
rect -45 3480 -30 3585
rect -80 3465 -30 3480
rect 20 3585 70 3600
rect 20 3480 35 3585
rect 55 3480 70 3585
rect 20 3465 70 3480
rect 120 3585 170 3600
rect 120 3480 135 3585
rect 155 3480 170 3585
rect 120 3465 170 3480
rect 220 3585 270 3600
rect 220 3480 235 3585
rect 255 3480 270 3585
rect 220 3465 270 3480
rect 320 3585 370 3600
rect 320 3480 335 3585
rect 355 3480 370 3585
rect 320 3465 370 3480
rect -680 2800 -630 2815
rect -680 2530 -665 2800
rect -645 2530 -630 2800
rect -680 2515 -630 2530
rect -580 2800 -530 2815
rect -580 2530 -565 2800
rect -545 2530 -530 2800
rect -580 2515 -530 2530
rect -480 2800 -430 2815
rect -480 2530 -465 2800
rect -445 2530 -430 2800
rect -480 2515 -430 2530
rect -380 2800 -330 2815
rect -380 2530 -365 2800
rect -345 2530 -330 2800
rect -380 2515 -330 2530
rect -280 2800 -230 2815
rect -280 2530 -265 2800
rect -245 2530 -230 2800
rect -280 2515 -230 2530
rect -180 2800 -130 2815
rect -180 2530 -165 2800
rect -145 2530 -130 2800
rect -180 2515 -130 2530
rect -80 2800 -30 2815
rect -80 2530 -65 2800
rect -45 2530 -30 2800
rect -80 2515 -30 2530
rect 20 2800 70 2815
rect 20 2530 35 2800
rect 55 2530 70 2800
rect 20 2515 70 2530
rect 120 2800 170 2815
rect 120 2530 135 2800
rect 155 2530 170 2800
rect 120 2515 170 2530
rect 220 2800 270 2815
rect 220 2530 235 2800
rect 255 2530 270 2800
rect 220 2515 270 2530
rect 320 2800 370 2815
rect 320 2530 335 2800
rect 355 2530 370 2800
rect 320 2515 370 2530
rect -680 1850 -630 1865
rect -680 1280 -665 1850
rect -645 1280 -630 1850
rect -680 1265 -630 1280
rect -580 1850 -530 1865
rect -580 1280 -565 1850
rect -545 1280 -530 1850
rect -580 1265 -530 1280
rect -480 1850 -430 1865
rect -480 1280 -465 1850
rect -445 1280 -430 1850
rect -480 1265 -430 1280
rect -380 1850 -330 1865
rect -380 1280 -365 1850
rect -345 1280 -330 1850
rect -380 1265 -330 1280
rect -280 1850 -230 1865
rect -280 1280 -265 1850
rect -245 1280 -230 1850
rect -280 1265 -230 1280
rect -180 1850 -130 1865
rect -180 1280 -165 1850
rect -145 1280 -130 1850
rect -180 1265 -130 1280
rect -80 1850 -30 1865
rect -80 1280 -65 1850
rect -45 1280 -30 1850
rect -80 1265 -30 1280
rect 20 1850 70 1865
rect 20 1280 35 1850
rect 55 1280 70 1850
rect 20 1265 70 1280
rect 120 1850 170 1865
rect 120 1280 135 1850
rect 155 1280 170 1850
rect 120 1265 170 1280
rect 220 1850 270 1865
rect 220 1280 235 1850
rect 255 1280 270 1850
rect 220 1265 270 1280
rect 320 1850 370 1865
rect 320 1280 335 1850
rect 355 1280 370 1850
rect 320 1265 370 1280
<< ndiffc >>
rect -665 30 -645 600
rect -565 30 -545 600
rect -465 30 -445 600
rect -365 30 -345 600
rect -265 30 -245 600
rect -165 30 -145 600
rect -65 30 -45 600
rect 35 30 55 600
rect 135 30 155 600
rect 235 30 255 600
rect 335 30 355 600
<< pdiffc >>
rect -665 3480 -645 3585
rect -565 3480 -545 3585
rect -465 3480 -445 3585
rect -365 3480 -345 3585
rect -265 3480 -245 3585
rect -165 3480 -145 3585
rect -65 3480 -45 3585
rect 35 3480 55 3585
rect 135 3480 155 3585
rect 235 3480 255 3585
rect 335 3480 355 3585
rect -665 2530 -645 2800
rect -565 2530 -545 2800
rect -465 2530 -445 2800
rect -365 2530 -345 2800
rect -265 2530 -245 2800
rect -165 2530 -145 2800
rect -65 2530 -45 2800
rect 35 2530 55 2800
rect 135 2530 155 2800
rect 235 2530 255 2800
rect 335 2530 355 2800
rect -665 1280 -645 1850
rect -565 1280 -545 1850
rect -465 1280 -445 1850
rect -365 1280 -345 1850
rect -265 1280 -245 1850
rect -165 1280 -145 1850
rect -65 1280 -45 1850
rect 35 1280 55 1850
rect 135 1280 155 1850
rect 235 1280 255 1850
rect 335 1280 355 1850
<< psubdiff >>
rect -730 600 -680 615
rect -730 30 -715 600
rect -695 30 -680 600
rect -730 15 -680 30
rect 370 600 420 615
rect 370 30 385 600
rect 405 30 420 600
rect 370 15 420 30
<< nsubdiff >>
rect -730 3585 -680 3600
rect -730 3480 -715 3585
rect -695 3480 -680 3585
rect -730 3465 -680 3480
rect 370 3585 420 3600
rect 370 3480 385 3585
rect 405 3480 420 3585
rect 370 3465 420 3480
rect -730 2800 -680 2815
rect -730 2530 -715 2800
rect -695 2530 -680 2800
rect -730 2515 -680 2530
rect 370 2800 420 2815
rect 370 2530 385 2800
rect 405 2530 420 2800
rect 370 2515 420 2530
rect -730 1850 -680 1865
rect -730 1280 -715 1850
rect -695 1280 -680 1850
rect -730 1265 -680 1280
rect 370 1850 420 1865
rect 370 1280 385 1850
rect 405 1280 420 1850
rect 370 1265 420 1280
<< psubdiffcont >>
rect -715 30 -695 600
rect 385 30 405 600
<< nsubdiffcont >>
rect -715 3480 -695 3585
rect 385 3480 405 3585
rect -715 2530 -695 2800
rect 385 2530 405 2800
rect -715 1280 -695 1850
rect 385 1280 405 1850
<< poly >>
rect -630 3600 -580 3615
rect -530 3600 -480 3615
rect -430 3600 -380 3615
rect -330 3600 -280 3615
rect -230 3600 -180 3615
rect -130 3600 -80 3615
rect -30 3600 20 3615
rect 70 3600 120 3615
rect 170 3600 220 3615
rect 270 3600 320 3615
rect -630 3450 -580 3465
rect -530 3450 -480 3465
rect -430 3450 -380 3465
rect -330 3450 -280 3465
rect -230 3450 -180 3465
rect -130 3450 -80 3465
rect -30 3450 20 3465
rect 70 3450 120 3465
rect 170 3450 220 3465
rect 270 3450 320 3465
rect -630 2815 -580 2830
rect -530 2815 -480 2830
rect -430 2815 -380 2830
rect -330 2815 -280 2830
rect -230 2815 -180 2830
rect -130 2815 -80 2830
rect -30 2815 20 2830
rect 70 2815 120 2830
rect 170 2815 220 2830
rect 270 2815 320 2830
rect -630 2500 -580 2515
rect -530 2500 -480 2515
rect -430 2500 -380 2515
rect -330 2500 -280 2515
rect -230 2500 -180 2515
rect -130 2500 -80 2515
rect -30 2500 20 2515
rect 70 2500 120 2515
rect 170 2500 220 2515
rect 270 2500 320 2515
rect -630 1865 -580 1880
rect -530 1865 -480 1880
rect -430 1865 -380 1880
rect -330 1865 -280 1880
rect -230 1865 -180 1880
rect -130 1865 -80 1880
rect -30 1865 20 1880
rect 70 1865 120 1880
rect 170 1865 220 1880
rect 270 1865 320 1880
rect -630 1250 -580 1265
rect -530 1250 -480 1265
rect -430 1250 -380 1265
rect -330 1250 -280 1265
rect -230 1250 -180 1265
rect -130 1250 -80 1265
rect -30 1250 20 1265
rect 70 1250 120 1265
rect 170 1250 220 1265
rect 270 1250 320 1265
rect -630 615 -580 630
rect -530 615 -480 630
rect -430 615 -380 630
rect -330 615 -280 630
rect -230 615 -180 630
rect -130 615 -80 630
rect -30 615 20 630
rect 70 615 120 630
rect 170 615 220 630
rect 270 615 320 630
rect -630 0 -580 15
rect -530 0 -480 15
rect -430 0 -380 15
rect -330 0 -280 15
rect -230 0 -180 15
rect -130 0 -80 15
rect -30 0 20 15
rect 70 0 120 15
rect 170 0 220 15
rect 270 0 320 15
<< locali >>
rect -725 3585 -635 3595
rect -725 3480 -715 3585
rect -695 3480 -665 3585
rect -645 3480 -635 3585
rect -725 3470 -635 3480
rect -575 3585 -535 3595
rect -575 3480 -565 3585
rect -545 3480 -535 3585
rect -575 3470 -535 3480
rect -475 3585 -435 3595
rect -475 3480 -465 3585
rect -445 3480 -435 3585
rect -475 3470 -435 3480
rect -375 3585 -335 3595
rect -375 3480 -365 3585
rect -345 3480 -335 3585
rect -375 3470 -335 3480
rect -275 3585 -235 3595
rect -275 3480 -265 3585
rect -245 3480 -235 3585
rect -275 3470 -235 3480
rect -175 3585 -135 3595
rect -175 3480 -165 3585
rect -145 3480 -135 3585
rect -175 3470 -135 3480
rect -75 3585 -35 3595
rect -75 3480 -65 3585
rect -45 3480 -35 3585
rect -75 3470 -35 3480
rect 25 3585 65 3595
rect 25 3480 35 3585
rect 55 3480 65 3585
rect 25 3470 65 3480
rect 125 3585 165 3595
rect 125 3480 135 3585
rect 155 3480 165 3585
rect 125 3470 165 3480
rect 225 3585 265 3595
rect 225 3480 235 3585
rect 255 3480 265 3585
rect 225 3470 265 3480
rect 325 3585 415 3595
rect 325 3480 335 3585
rect 355 3480 385 3585
rect 405 3480 415 3585
rect 325 3470 415 3480
rect -725 2800 -635 2810
rect -725 2530 -715 2800
rect -695 2530 -665 2800
rect -645 2530 -635 2800
rect -725 2520 -635 2530
rect -575 2800 -535 2810
rect -575 2530 -565 2800
rect -545 2530 -535 2800
rect -575 2520 -535 2530
rect -475 2800 -435 2810
rect -475 2530 -465 2800
rect -445 2530 -435 2800
rect -475 2520 -435 2530
rect -375 2800 -335 2810
rect -375 2530 -365 2800
rect -345 2530 -335 2800
rect -375 2520 -335 2530
rect -275 2800 -235 2810
rect -275 2530 -265 2800
rect -245 2530 -235 2800
rect -275 2520 -235 2530
rect -175 2800 -135 2810
rect -175 2530 -165 2800
rect -145 2530 -135 2800
rect -175 2520 -135 2530
rect -75 2800 -35 2810
rect -75 2530 -65 2800
rect -45 2530 -35 2800
rect -75 2520 -35 2530
rect 25 2800 65 2810
rect 25 2530 35 2800
rect 55 2530 65 2800
rect 25 2520 65 2530
rect 125 2800 165 2810
rect 125 2530 135 2800
rect 155 2530 165 2800
rect 125 2520 165 2530
rect 225 2800 265 2810
rect 225 2530 235 2800
rect 255 2530 265 2800
rect 225 2520 265 2530
rect 325 2800 415 2810
rect 325 2530 335 2800
rect 355 2530 385 2800
rect 405 2530 415 2800
rect 325 2520 415 2530
rect -725 1850 -635 1860
rect -725 1280 -715 1850
rect -695 1280 -665 1850
rect -645 1280 -635 1850
rect -725 1270 -635 1280
rect -575 1850 -535 1860
rect -575 1280 -565 1850
rect -545 1280 -535 1850
rect -575 1270 -535 1280
rect -475 1850 -435 1860
rect -475 1280 -465 1850
rect -445 1280 -435 1850
rect -475 1270 -435 1280
rect -375 1850 -335 1860
rect -375 1280 -365 1850
rect -345 1280 -335 1850
rect -375 1270 -335 1280
rect -275 1850 -235 1860
rect -275 1280 -265 1850
rect -245 1280 -235 1850
rect -275 1270 -235 1280
rect -175 1850 -135 1860
rect -175 1280 -165 1850
rect -145 1280 -135 1850
rect -175 1270 -135 1280
rect -75 1850 -35 1860
rect -75 1280 -65 1850
rect -45 1280 -35 1850
rect -75 1270 -35 1280
rect 25 1850 65 1860
rect 25 1280 35 1850
rect 55 1280 65 1850
rect 25 1270 65 1280
rect 125 1850 165 1860
rect 125 1280 135 1850
rect 155 1280 165 1850
rect 125 1270 165 1280
rect 225 1850 265 1860
rect 225 1280 235 1850
rect 255 1280 265 1850
rect 225 1270 265 1280
rect 325 1850 415 1860
rect 325 1280 335 1850
rect 355 1280 385 1850
rect 405 1280 415 1850
rect 325 1270 415 1280
rect -725 600 -635 610
rect -725 30 -715 600
rect -695 30 -665 600
rect -645 30 -635 600
rect -725 20 -635 30
rect -575 600 -535 610
rect -575 30 -565 600
rect -545 30 -535 600
rect -575 20 -535 30
rect -475 600 -435 610
rect -475 30 -465 600
rect -445 30 -435 600
rect -475 20 -435 30
rect -375 600 -335 610
rect -375 30 -365 600
rect -345 30 -335 600
rect -375 20 -335 30
rect -275 600 -235 610
rect -275 30 -265 600
rect -245 30 -235 600
rect -275 20 -235 30
rect -175 600 -135 610
rect -175 30 -165 600
rect -145 30 -135 600
rect -175 20 -135 30
rect -75 600 -35 610
rect -75 30 -65 600
rect -45 30 -35 600
rect -75 20 -35 30
rect 25 600 65 610
rect 25 30 35 600
rect 55 30 65 600
rect 25 20 65 30
rect 125 600 165 610
rect 125 30 135 600
rect 155 30 165 600
rect 125 20 165 30
rect 225 600 265 610
rect 225 30 235 600
rect 255 30 265 600
rect 225 20 265 30
rect 325 600 415 610
rect 325 30 335 600
rect 355 30 385 600
rect 405 30 415 600
rect 325 20 415 30
<< end >>
