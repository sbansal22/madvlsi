magic
tech sky130A
timestamp 1615885406
<< nwell >>
rect -750 1245 440 2855
<< nmos >>
rect -630 320 -580 920
rect -530 320 -480 920
rect -430 320 -380 920
rect -330 320 -280 920
rect -230 320 -180 920
rect -130 320 -80 920
rect -30 320 20 920
rect 70 320 120 920
rect 170 320 220 920
rect 270 320 320 920
<< pmos >>
rect -630 2700 -580 2835
rect -530 2700 -480 2835
rect -430 2700 -380 2835
rect -330 2700 -280 2835
rect -230 2700 -180 2835
rect -130 2700 -80 2835
rect -30 2700 20 2835
rect 70 2700 120 2835
rect 170 2700 220 2835
rect 270 2700 320 2835
rect -630 2145 -580 2445
rect -530 2145 -480 2445
rect -430 2145 -380 2445
rect -330 2145 -280 2445
rect -230 2145 -180 2445
rect -130 2145 -80 2445
rect -30 2145 20 2445
rect 70 2145 120 2445
rect 170 2145 220 2445
rect 270 2145 320 2445
rect -630 1265 -580 1865
rect -530 1265 -480 1865
rect -430 1265 -380 1865
rect -330 1265 -280 1865
rect -230 1265 -180 1865
rect -130 1265 -80 1865
rect -30 1265 20 1865
rect 70 1265 120 1865
rect 170 1265 220 1865
rect 270 1265 320 1865
<< ndiff >>
rect -680 905 -630 920
rect -680 335 -665 905
rect -645 335 -630 905
rect -680 320 -630 335
rect -580 905 -530 920
rect -580 335 -565 905
rect -545 335 -530 905
rect -580 320 -530 335
rect -480 905 -430 920
rect -480 335 -465 905
rect -445 335 -430 905
rect -480 320 -430 335
rect -380 905 -330 920
rect -380 335 -365 905
rect -345 335 -330 905
rect -380 320 -330 335
rect -280 905 -230 920
rect -280 335 -265 905
rect -245 335 -230 905
rect -280 320 -230 335
rect -180 905 -130 920
rect -180 335 -165 905
rect -145 335 -130 905
rect -180 320 -130 335
rect -80 905 -30 920
rect -80 335 -65 905
rect -45 335 -30 905
rect -80 320 -30 335
rect 20 905 70 920
rect 20 335 35 905
rect 55 335 70 905
rect 20 320 70 335
rect 120 905 170 920
rect 120 335 135 905
rect 155 335 170 905
rect 120 320 170 335
rect 220 905 270 920
rect 220 335 235 905
rect 255 335 270 905
rect 220 320 270 335
rect 320 905 370 920
rect 320 335 335 905
rect 355 335 370 905
rect 320 320 370 335
<< pdiff >>
rect -680 2820 -630 2835
rect -680 2715 -665 2820
rect -645 2715 -630 2820
rect -680 2700 -630 2715
rect -580 2820 -530 2835
rect -580 2715 -565 2820
rect -545 2715 -530 2820
rect -580 2700 -530 2715
rect -480 2820 -430 2835
rect -480 2715 -465 2820
rect -445 2715 -430 2820
rect -480 2700 -430 2715
rect -380 2820 -330 2835
rect -380 2715 -365 2820
rect -345 2715 -330 2820
rect -380 2700 -330 2715
rect -280 2820 -230 2835
rect -280 2715 -265 2820
rect -245 2715 -230 2820
rect -280 2700 -230 2715
rect -180 2820 -130 2835
rect -180 2715 -165 2820
rect -145 2715 -130 2820
rect -180 2700 -130 2715
rect -80 2820 -30 2835
rect -80 2715 -65 2820
rect -45 2715 -30 2820
rect -80 2700 -30 2715
rect 20 2820 70 2835
rect 20 2715 35 2820
rect 55 2715 70 2820
rect 20 2700 70 2715
rect 120 2820 170 2835
rect 120 2715 135 2820
rect 155 2715 170 2820
rect 120 2700 170 2715
rect 220 2820 270 2835
rect 220 2715 235 2820
rect 255 2715 270 2820
rect 220 2700 270 2715
rect 320 2820 370 2835
rect 320 2715 335 2820
rect 355 2715 370 2820
rect 320 2700 370 2715
rect -680 2430 -630 2445
rect -680 2160 -665 2430
rect -645 2160 -630 2430
rect -680 2145 -630 2160
rect -580 2430 -530 2445
rect -580 2160 -565 2430
rect -545 2160 -530 2430
rect -580 2145 -530 2160
rect -480 2430 -430 2445
rect -480 2160 -465 2430
rect -445 2160 -430 2430
rect -480 2145 -430 2160
rect -380 2430 -330 2445
rect -380 2160 -365 2430
rect -345 2160 -330 2430
rect -380 2145 -330 2160
rect -280 2430 -230 2445
rect -280 2160 -265 2430
rect -245 2160 -230 2430
rect -280 2145 -230 2160
rect -180 2430 -130 2445
rect -180 2160 -165 2430
rect -145 2160 -130 2430
rect -180 2145 -130 2160
rect -80 2430 -30 2445
rect -80 2160 -65 2430
rect -45 2160 -30 2430
rect -80 2145 -30 2160
rect 20 2430 70 2445
rect 20 2160 35 2430
rect 55 2160 70 2430
rect 20 2145 70 2160
rect 120 2430 170 2445
rect 120 2160 135 2430
rect 155 2160 170 2430
rect 120 2145 170 2160
rect 220 2430 270 2445
rect 220 2160 235 2430
rect 255 2160 270 2430
rect 220 2145 270 2160
rect 320 2430 370 2445
rect 320 2160 335 2430
rect 355 2160 370 2430
rect 320 2145 370 2160
rect -680 1850 -630 1865
rect -680 1280 -665 1850
rect -645 1280 -630 1850
rect -680 1265 -630 1280
rect -580 1850 -530 1865
rect -580 1280 -565 1850
rect -545 1280 -530 1850
rect -580 1265 -530 1280
rect -480 1850 -430 1865
rect -480 1280 -465 1850
rect -445 1280 -430 1850
rect -480 1265 -430 1280
rect -380 1850 -330 1865
rect -380 1280 -365 1850
rect -345 1280 -330 1850
rect -380 1265 -330 1280
rect -280 1850 -230 1865
rect -280 1280 -265 1850
rect -245 1280 -230 1850
rect -280 1265 -230 1280
rect -180 1850 -130 1865
rect -180 1280 -165 1850
rect -145 1280 -130 1850
rect -180 1265 -130 1280
rect -80 1850 -30 1865
rect -80 1280 -65 1850
rect -45 1280 -30 1850
rect -80 1265 -30 1280
rect 20 1850 70 1865
rect 20 1280 35 1850
rect 55 1280 70 1850
rect 20 1265 70 1280
rect 120 1850 170 1865
rect 120 1280 135 1850
rect 155 1280 170 1850
rect 120 1265 170 1280
rect 220 1850 270 1865
rect 220 1280 235 1850
rect 255 1280 270 1850
rect 220 1265 270 1280
rect 320 1850 370 1865
rect 320 1280 335 1850
rect 355 1280 370 1850
rect 320 1265 370 1280
<< ndiffc >>
rect -665 335 -645 905
rect -565 335 -545 905
rect -465 335 -445 905
rect -365 335 -345 905
rect -265 335 -245 905
rect -165 335 -145 905
rect -65 335 -45 905
rect 35 335 55 905
rect 135 335 155 905
rect 235 335 255 905
rect 335 335 355 905
<< pdiffc >>
rect -665 2715 -645 2820
rect -565 2715 -545 2820
rect -465 2715 -445 2820
rect -365 2715 -345 2820
rect -265 2715 -245 2820
rect -165 2715 -145 2820
rect -65 2715 -45 2820
rect 35 2715 55 2820
rect 135 2715 155 2820
rect 235 2715 255 2820
rect 335 2715 355 2820
rect -665 2160 -645 2430
rect -565 2160 -545 2430
rect -465 2160 -445 2430
rect -365 2160 -345 2430
rect -265 2160 -245 2430
rect -165 2160 -145 2430
rect -65 2160 -45 2430
rect 35 2160 55 2430
rect 135 2160 155 2430
rect 235 2160 255 2430
rect 335 2160 355 2430
rect -665 1280 -645 1850
rect -565 1280 -545 1850
rect -465 1280 -445 1850
rect -365 1280 -345 1850
rect -265 1280 -245 1850
rect -165 1280 -145 1850
rect -65 1280 -45 1850
rect 35 1280 55 1850
rect 135 1280 155 1850
rect 235 1280 255 1850
rect 335 1280 355 1850
<< psubdiff >>
rect -730 905 -680 920
rect -730 335 -715 905
rect -695 335 -680 905
rect -730 320 -680 335
rect 370 905 420 920
rect 370 335 385 905
rect 405 335 420 905
rect 370 320 420 335
<< nsubdiff >>
rect -730 2820 -680 2835
rect -730 2715 -715 2820
rect -695 2715 -680 2820
rect -730 2700 -680 2715
rect 370 2820 420 2835
rect 370 2715 385 2820
rect 405 2715 420 2820
rect 370 2700 420 2715
rect -730 2430 -680 2445
rect -730 2160 -715 2430
rect -695 2160 -680 2430
rect -730 2145 -680 2160
rect 370 2430 420 2445
rect 370 2160 385 2430
rect 405 2160 420 2430
rect 370 2145 420 2160
rect -730 1850 -680 1865
rect -730 1280 -715 1850
rect -695 1280 -680 1850
rect -730 1265 -680 1280
rect 370 1850 420 1865
rect 370 1280 385 1850
rect 405 1280 420 1850
rect 370 1265 420 1280
<< psubdiffcont >>
rect -715 335 -695 905
rect 385 335 405 905
<< nsubdiffcont >>
rect -715 2715 -695 2820
rect 385 2715 405 2820
rect -715 2160 -695 2430
rect 385 2160 405 2430
rect -715 1280 -695 1850
rect 385 1280 405 1850
<< poly >>
rect -630 2835 -580 2850
rect -530 2835 -480 2850
rect -430 2835 -380 2850
rect -330 2835 -280 2850
rect -230 2835 -180 2850
rect -130 2835 -80 2850
rect -30 2835 20 2850
rect 70 2835 120 2850
rect 170 2835 220 2850
rect 270 2835 320 2850
rect -630 2685 -580 2700
rect -530 2685 -480 2700
rect -430 2685 -380 2700
rect -330 2685 -280 2700
rect -230 2685 -180 2700
rect -130 2685 -80 2700
rect -30 2685 20 2700
rect 70 2685 120 2700
rect 170 2685 220 2700
rect -675 2675 -580 2685
rect -675 2655 -665 2675
rect -645 2670 -580 2675
rect -555 2670 220 2685
rect 270 2685 320 2700
rect 270 2675 365 2685
rect 270 2670 335 2675
rect -645 2655 -635 2670
rect -675 2645 -635 2655
rect -555 2620 -540 2670
rect 325 2655 335 2670
rect 355 2655 365 2675
rect 325 2645 365 2655
rect -730 2610 -540 2620
rect -730 2590 -720 2610
rect -700 2605 -540 2610
rect -700 2590 -690 2605
rect -730 2580 -690 2590
rect -730 2545 -380 2555
rect -730 2525 -720 2545
rect -700 2540 -380 2545
rect -700 2525 -690 2540
rect -730 2515 -690 2525
rect -430 2500 -380 2540
rect -675 2490 -635 2500
rect -675 2470 -665 2490
rect -645 2475 -635 2490
rect -430 2485 120 2500
rect -645 2470 -580 2475
rect -675 2460 -580 2470
rect -630 2445 -580 2460
rect -530 2445 -480 2460
rect -430 2445 -380 2485
rect -330 2445 -280 2485
rect -230 2445 -180 2460
rect -130 2445 -80 2460
rect -30 2445 20 2485
rect 70 2445 120 2485
rect 325 2490 365 2500
rect 325 2475 335 2490
rect 270 2470 335 2475
rect 355 2470 365 2490
rect 270 2460 365 2470
rect 170 2445 220 2460
rect 270 2445 320 2460
rect -630 2130 -580 2145
rect -530 2105 -480 2145
rect -430 2130 -380 2145
rect -330 2130 -280 2145
rect -230 2105 -180 2145
rect -130 2105 -80 2145
rect -30 2130 20 2145
rect 70 2130 120 2145
rect 170 2105 220 2145
rect 270 2130 320 2145
rect -730 2095 220 2105
rect -730 2075 -720 2095
rect -700 2090 220 2095
rect -700 2075 -690 2090
rect -730 2065 -690 2075
rect -375 2055 65 2065
rect -375 2035 -365 2055
rect -345 2050 35 2055
rect -345 2035 -335 2050
rect -375 2025 -335 2035
rect 25 2035 35 2050
rect 55 2035 65 2055
rect 25 2025 65 2035
rect -575 2015 -535 2025
rect -575 1995 -565 2015
rect -545 1995 -535 2015
rect -575 1985 -535 1995
rect -730 1970 -620 1980
rect -730 1950 -720 1970
rect -700 1965 -620 1970
rect -700 1950 -690 1965
rect -730 1940 -690 1950
rect -635 1960 -620 1965
rect -635 1945 220 1960
rect -675 1910 -635 1920
rect -675 1890 -665 1910
rect -645 1895 -635 1910
rect -645 1890 -580 1895
rect -675 1880 -580 1890
rect -630 1865 -580 1880
rect -530 1865 -480 1945
rect -430 1865 -380 1880
rect -330 1865 -280 1880
rect -230 1865 -180 1945
rect -130 1865 -80 1945
rect -30 1865 20 1880
rect 70 1865 120 1880
rect 170 1865 220 1945
rect 325 1910 365 1920
rect 325 1895 335 1910
rect 270 1890 335 1895
rect 355 1890 365 1910
rect 270 1880 365 1890
rect 270 1865 320 1880
rect -630 1250 -580 1265
rect -530 1250 -480 1265
rect -430 1225 -380 1265
rect -330 1225 -280 1265
rect -230 1250 -180 1265
rect -130 1250 -80 1265
rect -30 1225 20 1265
rect 70 1225 120 1265
rect 170 1250 220 1265
rect 270 1250 320 1265
rect -430 1215 120 1225
rect -430 1210 -165 1215
rect -430 1120 -415 1210
rect -175 1195 -165 1210
rect -145 1210 120 1215
rect -145 1195 -135 1210
rect -175 1185 -135 1195
rect -575 1110 -415 1120
rect -575 1090 -565 1110
rect -545 1105 -415 1110
rect 105 1120 120 1210
rect 105 1110 265 1120
rect 105 1105 235 1110
rect -545 1090 -535 1105
rect -575 1080 -535 1090
rect 225 1090 235 1105
rect 255 1090 265 1110
rect 225 1080 265 1090
rect -725 1030 -685 1040
rect -725 1010 -715 1030
rect -695 1015 -685 1030
rect -695 1010 -415 1015
rect -725 1000 -415 1010
rect -430 975 -415 1000
rect -675 965 -635 975
rect -675 945 -665 965
rect -645 950 -635 965
rect -430 960 120 975
rect -645 945 -580 950
rect -675 935 -580 945
rect -630 920 -580 935
rect -530 920 -480 935
rect -430 920 -380 960
rect -330 920 -280 960
rect -230 920 -180 935
rect -130 920 -80 935
rect -30 920 20 960
rect 70 920 120 960
rect 325 965 365 975
rect 325 950 335 965
rect 270 945 335 950
rect 355 945 365 965
rect 270 935 365 945
rect 170 920 220 935
rect 270 920 320 935
rect -630 305 -580 320
rect -700 295 -660 305
rect -700 275 -690 295
rect -670 280 -660 295
rect -530 280 -480 320
rect -430 305 -380 320
rect -330 305 -280 320
rect -230 280 -180 320
rect -130 280 -80 320
rect -30 305 20 320
rect 70 305 120 320
rect 170 280 220 320
rect 270 305 320 320
rect -670 275 220 280
rect -700 265 220 275
<< polycont >>
rect -665 2655 -645 2675
rect 335 2655 355 2675
rect -720 2590 -700 2610
rect -720 2525 -700 2545
rect -665 2470 -645 2490
rect 335 2470 355 2490
rect -720 2075 -700 2095
rect -365 2035 -345 2055
rect 35 2035 55 2055
rect -565 1995 -545 2015
rect -720 1950 -700 1970
rect -665 1890 -645 1910
rect 335 1890 355 1910
rect -165 1195 -145 1215
rect -565 1090 -545 1110
rect 235 1090 255 1110
rect -715 1010 -695 1030
rect -665 945 -645 965
rect 335 945 355 965
rect -690 275 -670 295
<< locali >>
rect -725 2820 -635 2830
rect -725 2715 -715 2820
rect -695 2715 -665 2820
rect -645 2715 -635 2820
rect -725 2705 -635 2715
rect -575 2820 -535 2830
rect -575 2715 -565 2820
rect -545 2715 -535 2820
rect -575 2705 -535 2715
rect -475 2820 -435 2830
rect -475 2715 -465 2820
rect -445 2715 -435 2820
rect -675 2675 -635 2705
rect -675 2655 -665 2675
rect -645 2655 -635 2675
rect -675 2645 -635 2655
rect -475 2675 -435 2715
rect -375 2820 -335 2830
rect -375 2715 -365 2820
rect -345 2715 -335 2820
rect -375 2705 -335 2715
rect -275 2820 -235 2830
rect -275 2715 -265 2820
rect -245 2715 -235 2820
rect -275 2675 -235 2715
rect -175 2820 -135 2830
rect -175 2715 -165 2820
rect -145 2715 -135 2820
rect -175 2705 -135 2715
rect -75 2820 -35 2830
rect -75 2715 -65 2820
rect -45 2715 -35 2820
rect -75 2675 -35 2715
rect 25 2820 65 2830
rect 25 2715 35 2820
rect 55 2715 65 2820
rect 25 2705 65 2715
rect 125 2820 165 2830
rect 125 2715 135 2820
rect 155 2715 165 2820
rect 125 2675 165 2715
rect 225 2820 265 2830
rect 225 2715 235 2820
rect 255 2715 265 2820
rect 225 2705 265 2715
rect 325 2820 415 2830
rect 325 2715 335 2820
rect 355 2715 385 2820
rect 405 2715 415 2820
rect 325 2705 415 2715
rect -475 2655 165 2675
rect -750 2610 -690 2620
rect -750 2600 -720 2610
rect -730 2590 -720 2600
rect -700 2590 -690 2610
rect -730 2580 -690 2590
rect -750 2545 -690 2555
rect -750 2535 -720 2545
rect -730 2525 -720 2535
rect -700 2525 -690 2545
rect -730 2515 -690 2525
rect -675 2490 -635 2500
rect -675 2470 -665 2490
rect -645 2470 -635 2490
rect -675 2440 -635 2470
rect -725 2430 -635 2440
rect -725 2160 -715 2430
rect -695 2160 -665 2430
rect -645 2160 -635 2430
rect -725 2150 -635 2160
rect -575 2430 -535 2440
rect -575 2160 -565 2430
rect -545 2160 -535 2430
rect -750 2095 -690 2105
rect -750 2085 -720 2095
rect -730 2075 -720 2085
rect -700 2075 -690 2095
rect -730 2065 -690 2075
rect -575 2015 -535 2160
rect -475 2430 -435 2655
rect -475 2160 -465 2430
rect -445 2160 -435 2430
rect -475 2150 -435 2160
rect -375 2430 -335 2440
rect -375 2160 -365 2430
rect -345 2160 -335 2430
rect -375 2065 -335 2160
rect -275 2430 -235 2655
rect -275 2160 -265 2430
rect -245 2160 -235 2430
rect -275 2150 -235 2160
rect -175 2430 -135 2440
rect -175 2160 -165 2430
rect -145 2160 -135 2430
rect -440 2055 -335 2065
rect -440 2035 -430 2055
rect -410 2045 -365 2055
rect -410 2035 -400 2045
rect -440 2025 -400 2035
rect -375 2035 -365 2045
rect -345 2035 -335 2055
rect -375 2025 -335 2035
rect -575 1995 -565 2015
rect -545 2005 -535 2015
rect -175 2015 -135 2160
rect -75 2430 -35 2655
rect -75 2160 -65 2430
rect -45 2160 -35 2430
rect -75 2150 -35 2160
rect 25 2430 65 2440
rect 25 2160 35 2430
rect 55 2160 65 2430
rect 25 2055 65 2160
rect 125 2430 165 2655
rect 325 2675 365 2705
rect 325 2655 335 2675
rect 355 2655 365 2675
rect 325 2645 365 2655
rect 325 2490 365 2500
rect 325 2470 335 2490
rect 355 2470 365 2490
rect 325 2440 365 2470
rect 125 2160 135 2430
rect 155 2160 165 2430
rect 125 2150 165 2160
rect 225 2430 265 2440
rect 225 2160 235 2430
rect 255 2160 265 2430
rect 25 2035 35 2055
rect 55 2035 65 2055
rect 25 2025 65 2035
rect -175 2005 -165 2015
rect -545 1995 -165 2005
rect -145 2005 -135 2015
rect 225 2005 265 2160
rect 325 2430 415 2440
rect 325 2160 335 2430
rect 355 2160 385 2430
rect 405 2160 415 2430
rect 325 2150 415 2160
rect -145 1995 265 2005
rect -575 1985 265 1995
rect -750 1970 -690 1980
rect -750 1955 -720 1970
rect -730 1950 -720 1955
rect -700 1950 -690 1970
rect -730 1940 -690 1950
rect -475 1920 165 1940
rect -675 1910 -635 1920
rect -675 1890 -665 1910
rect -645 1890 -635 1910
rect -675 1860 -635 1890
rect -725 1850 -635 1860
rect -725 1280 -715 1850
rect -695 1280 -665 1850
rect -645 1280 -635 1850
rect -725 1270 -635 1280
rect -575 1850 -535 1860
rect -575 1280 -565 1850
rect -545 1280 -535 1850
rect -575 1165 -535 1280
rect -475 1850 -435 1920
rect -275 1880 -35 1900
rect -475 1280 -465 1850
rect -445 1280 -435 1850
rect -475 1270 -435 1280
rect -375 1850 -335 1860
rect -375 1280 -365 1850
rect -345 1280 -335 1850
rect -375 1270 -335 1280
rect -275 1850 -235 1880
rect -275 1280 -265 1850
rect -245 1280 -235 1850
rect -275 1270 -235 1280
rect -175 1850 -135 1860
rect -175 1280 -165 1850
rect -145 1280 -135 1850
rect -175 1215 -135 1280
rect -75 1850 -35 1880
rect -75 1280 -65 1850
rect -45 1280 -35 1850
rect -75 1270 -35 1280
rect 25 1850 65 1860
rect 25 1280 35 1850
rect 55 1280 65 1850
rect 25 1270 65 1280
rect 125 1850 165 1920
rect 325 1910 365 1920
rect 325 1890 335 1910
rect 355 1890 365 1910
rect 325 1865 365 1890
rect 325 1860 370 1865
rect 125 1280 135 1850
rect 155 1280 165 1850
rect 125 1270 165 1280
rect 225 1850 265 1860
rect 225 1280 235 1850
rect 255 1280 265 1850
rect -175 1195 -165 1215
rect -145 1195 -135 1215
rect -175 1185 -135 1195
rect 225 1165 265 1280
rect 325 1850 415 1860
rect 325 1280 335 1850
rect 355 1280 385 1850
rect 405 1280 415 1850
rect 325 1270 415 1280
rect -575 1145 440 1165
rect -575 1110 -535 1120
rect -575 1090 -565 1110
rect -545 1090 -535 1110
rect -725 1030 -685 1040
rect -725 1020 -715 1030
rect -730 1010 -715 1020
rect -695 1010 -685 1030
rect -730 1000 -685 1010
rect -675 965 -635 975
rect -675 945 -665 965
rect -645 945 -635 965
rect -675 920 -635 945
rect -680 915 -635 920
rect -725 905 -635 915
rect -725 335 -715 905
rect -695 335 -665 905
rect -645 335 -635 905
rect -725 325 -635 335
rect -575 905 -535 1090
rect -575 335 -565 905
rect -545 335 -535 905
rect -575 325 -535 335
rect -475 1070 -435 1080
rect -475 1050 -465 1070
rect -445 1050 -435 1070
rect -475 905 -435 1050
rect -475 335 -465 905
rect -445 335 -435 905
rect -700 295 -660 305
rect -700 285 -690 295
rect -730 275 -690 285
rect -670 275 -660 295
rect -730 265 -660 275
rect -475 265 -435 335
rect -375 905 -335 915
rect -375 335 -365 905
rect -345 335 -335 905
rect -375 325 -335 335
rect -275 905 -235 915
rect -275 335 -265 905
rect -245 335 -235 905
rect -275 305 -235 335
rect -175 905 -135 1145
rect 225 1110 265 1120
rect 225 1090 235 1110
rect 255 1090 265 1110
rect -175 335 -165 905
rect -145 335 -135 905
rect -175 325 -135 335
rect -75 1030 -35 1040
rect -75 1010 -65 1030
rect -45 1010 -35 1030
rect -75 905 -35 1010
rect -75 335 -65 905
rect -45 335 -35 905
rect -75 305 -35 335
rect 25 905 65 915
rect 25 335 35 905
rect 55 335 65 905
rect 25 325 65 335
rect 125 905 165 915
rect 125 335 135 905
rect 155 335 165 905
rect -275 285 -35 305
rect 125 265 165 335
rect 225 905 265 1090
rect 225 335 235 905
rect 255 335 265 905
rect 225 325 265 335
rect 325 965 365 975
rect 325 945 335 965
rect 355 945 365 965
rect 325 915 365 945
rect 325 905 415 915
rect 325 335 335 905
rect 355 335 385 905
rect 405 335 415 905
rect 325 325 415 335
rect -475 245 165 265
<< viali >>
rect -715 2715 -695 2820
rect -665 2715 -645 2820
rect -565 2715 -545 2820
rect -365 2715 -345 2820
rect -165 2715 -145 2820
rect 35 2715 55 2820
rect 235 2715 255 2820
rect 335 2715 355 2820
rect 385 2715 405 2820
rect -430 2035 -410 2055
rect -165 1995 -145 2015
rect -715 1280 -695 1850
rect -665 1280 -645 1850
rect -365 1280 -345 1850
rect 35 1280 55 1850
rect 335 1280 355 1850
rect 385 1280 405 1850
rect -715 335 -695 905
rect -665 335 -645 905
rect -465 1050 -445 1070
rect -365 335 -345 905
rect -65 1010 -45 1030
rect 35 335 55 905
rect 335 335 355 905
rect 385 335 405 905
<< metal1 >>
rect -730 2820 420 2830
rect -730 2715 -715 2820
rect -695 2715 -665 2820
rect -645 2715 -565 2820
rect -545 2715 -365 2820
rect -345 2715 -165 2820
rect -145 2715 35 2820
rect 55 2715 235 2820
rect 255 2715 335 2820
rect 355 2715 385 2820
rect 405 2715 420 2820
rect -730 2150 420 2715
rect -730 1860 -635 2150
rect -440 2055 -400 2065
rect -440 2035 -430 2055
rect -410 2035 -400 2055
rect -440 1930 -400 2035
rect -175 2015 -135 2025
rect -175 1995 -165 2015
rect -145 1995 -135 2015
rect -175 1930 -135 1995
rect -440 1890 -235 1930
rect -175 1890 -35 1930
rect -730 1850 -335 1860
rect -730 1280 -715 1850
rect -695 1280 -665 1850
rect -645 1280 -365 1850
rect -345 1280 -335 1850
rect -730 1270 -335 1280
rect -275 1080 -235 1890
rect -475 1070 -235 1080
rect -475 1050 -465 1070
rect -445 1050 -235 1070
rect -475 1040 -235 1050
rect -75 1030 -35 1890
rect 325 1860 420 2150
rect 25 1850 420 1860
rect 25 1280 35 1850
rect 55 1280 335 1850
rect 355 1280 385 1850
rect 405 1280 420 1850
rect 25 1270 420 1280
rect -75 1010 -65 1030
rect -45 1010 -35 1030
rect -75 1000 -35 1010
rect -725 905 415 915
rect -725 335 -715 905
rect -695 335 -665 905
rect -645 335 -365 905
rect -345 335 35 905
rect 55 335 335 905
rect 355 335 385 905
rect 405 335 415 905
rect -725 325 415 335
<< end >>
